LVDS_TX_inst : LVDS_TX PORT MAP (
		pll_areset	 => pll_areset_sig,
		tx_in	 => tx_in_sig,
		tx_inclock	 => tx_inclock_sig,
		tx_out	 => tx_out_sig,
		tx_outclock	 => tx_outclock_sig
	);

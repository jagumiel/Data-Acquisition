LVDS_RX_inst : LVDS_RX PORT MAP (
		rx_in	 => rx_in_sig,
		rx_inclock	 => rx_inclock_sig,
		rx_out	 => rx_out_sig,
		rx_outclock	 => rx_outclock_sig
	);

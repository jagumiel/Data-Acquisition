library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use ieee.numeric_std.all;
--use ieee.numeric_std;


entity triangle is
	port (
		clk:		in	std_logic;
		amp:		in	std_logic_vector(32-1 downto 0);
		frq:		in	std_logic_vector(32-1 downto 0);
		pwm_ctrl:	out	std_logic_vector(32-1 downto 0)
	);
end triangle;

architecture Behavioral of triangle is

	type  SAMPLE_main is array (1 to 10000) of std_logic_vector(31 downto 0);--antes 1 to 100
	constant data : SAMPLE_main := (
		x"00000002",x"00000004",x"00000006",x"00000008",x"0000000a",x"0000000c",x"0000000e",x"00000010",
		x"00000012",x"00000014",x"00000016",x"00000018",x"0000001a",x"0000001c",x"0000001e",x"00000020",
		x"00000022",x"00000024",x"00000026",x"00000028",x"0000002a",x"0000002c",x"0000002e",x"00000030",
		x"00000032",x"00000034",x"00000036",x"00000038",x"0000003a",x"0000003c",x"0000003e",x"00000040",
		x"00000042",x"00000044",x"00000046",x"00000048",x"0000004a",x"0000004c",x"0000004e",x"00000050",
		x"00000052",x"00000054",x"00000056",x"00000058",x"0000005a",x"0000005c",x"0000005e",x"00000060",
		x"00000062",x"00000064",x"00000066",x"00000068",x"0000006a",x"0000006c",x"0000006e",x"00000070",
		x"00000072",x"00000074",x"00000076",x"00000078",x"0000007a",x"0000007c",x"0000007e",x"00000080",
		x"00000082",x"00000084",x"00000086",x"00000088",x"0000008a",x"0000008c",x"0000008e",x"00000090",
		x"00000092",x"00000094",x"00000096",x"00000098",x"0000009a",x"0000009c",x"0000009e",x"000000a0",
		x"000000a2",x"000000a4",x"000000a6",x"000000a8",x"000000aa",x"000000ac",x"000000ae",x"000000b0",
		x"000000b2",x"000000b4",x"000000b6",x"000000b8",x"000000ba",x"000000bc",x"000000be",x"000000c0",
		x"000000c2",x"000000c4",x"000000c6",x"000000c8",x"000000ca",x"000000cc",x"000000ce",x"000000d0",
		x"000000d2",x"000000d4",x"000000d6",x"000000d8",x"000000da",x"000000dc",x"000000de",x"000000e0",
		x"000000e2",x"000000e4",x"000000e6",x"000000e8",x"000000ea",x"000000ec",x"000000ee",x"000000f0",
		x"000000f2",x"000000f4",x"000000f6",x"000000f8",x"000000fa",x"000000fc",x"000000fe",x"00000100",
		x"00000102",x"00000104",x"00000106",x"00000108",x"0000010a",x"0000010c",x"0000010e",x"00000110",
		x"00000112",x"00000114",x"00000116",x"00000118",x"0000011a",x"0000011c",x"0000011e",x"00000120",
		x"00000122",x"00000124",x"00000126",x"00000128",x"0000012a",x"0000012c",x"0000012e",x"00000130",
		x"00000132",x"00000134",x"00000136",x"00000138",x"0000013a",x"0000013c",x"0000013e",x"00000140",
		x"00000142",x"00000144",x"00000146",x"00000148",x"0000014a",x"0000014c",x"0000014e",x"00000150",
		x"00000152",x"00000154",x"00000156",x"00000158",x"0000015a",x"0000015c",x"0000015e",x"00000160",
		x"00000162",x"00000164",x"00000166",x"00000168",x"0000016a",x"0000016c",x"0000016e",x"00000170",
		x"00000172",x"00000174",x"00000176",x"00000178",x"0000017a",x"0000017c",x"0000017e",x"00000180",
		x"00000182",x"00000184",x"00000186",x"00000188",x"0000018a",x"0000018c",x"0000018e",x"00000190",
		x"00000192",x"00000194",x"00000196",x"00000198",x"0000019a",x"0000019c",x"0000019e",x"000001a0",
		x"000001a2",x"000001a4",x"000001a6",x"000001a8",x"000001aa",x"000001ac",x"000001ae",x"000001b0",
		x"000001b2",x"000001b4",x"000001b6",x"000001b8",x"000001ba",x"000001bc",x"000001be",x"000001c0",
		x"000001c2",x"000001c4",x"000001c6",x"000001c8",x"000001ca",x"000001cc",x"000001ce",x"000001d0",
		x"000001d2",x"000001d4",x"000001d6",x"000001d8",x"000001da",x"000001dc",x"000001de",x"000001e0",
		x"000001e2",x"000001e4",x"000001e6",x"000001e8",x"000001ea",x"000001ec",x"000001ee",x"000001f0",
		x"000001f2",x"000001f4",x"000001f6",x"000001f8",x"000001fa",x"000001fc",x"000001fe",x"00000200",
		x"00000202",x"00000204",x"00000206",x"00000208",x"0000020a",x"0000020c",x"0000020e",x"00000210",
		x"00000212",x"00000214",x"00000216",x"00000218",x"0000021a",x"0000021c",x"0000021e",x"00000220",
		x"00000222",x"00000224",x"00000226",x"00000228",x"0000022a",x"0000022c",x"0000022e",x"00000230",
		x"00000232",x"00000234",x"00000236",x"00000238",x"0000023a",x"0000023c",x"0000023e",x"00000240",
		x"00000242",x"00000244",x"00000246",x"00000248",x"0000024a",x"0000024c",x"0000024e",x"00000250",
		x"00000252",x"00000254",x"00000256",x"00000258",x"0000025a",x"0000025c",x"0000025e",x"00000260",
		x"00000262",x"00000264",x"00000266",x"00000268",x"0000026a",x"0000026c",x"0000026e",x"00000270",
		x"00000272",x"00000274",x"00000276",x"00000278",x"0000027a",x"0000027c",x"0000027e",x"00000280",
		x"00000282",x"00000284",x"00000286",x"00000288",x"0000028a",x"0000028c",x"0000028e",x"00000290",
		x"00000292",x"00000294",x"00000296",x"00000298",x"0000029a",x"0000029c",x"0000029e",x"000002a0",
		x"000002a2",x"000002a4",x"000002a6",x"000002a8",x"000002aa",x"000002ac",x"000002ae",x"000002b0",
		x"000002b2",x"000002b4",x"000002b6",x"000002b8",x"000002ba",x"000002bc",x"000002be",x"000002c0",
		x"000002c2",x"000002c4",x"000002c6",x"000002c8",x"000002ca",x"000002cc",x"000002ce",x"000002d0",
		x"000002d2",x"000002d4",x"000002d6",x"000002d8",x"000002da",x"000002dc",x"000002de",x"000002e0",
		x"000002e2",x"000002e4",x"000002e6",x"000002e8",x"000002ea",x"000002ec",x"000002ee",x"000002f0",
		x"000002f2",x"000002f4",x"000002f6",x"000002f8",x"000002fa",x"000002fc",x"000002fe",x"00000300",
		x"00000302",x"00000304",x"00000306",x"00000308",x"0000030a",x"0000030c",x"0000030e",x"00000310",
		x"00000312",x"00000314",x"00000316",x"00000318",x"0000031a",x"0000031c",x"0000031e",x"00000320",
		x"00000322",x"00000324",x"00000326",x"00000328",x"0000032a",x"0000032c",x"0000032e",x"00000330",
		x"00000332",x"00000334",x"00000336",x"00000338",x"0000033a",x"0000033c",x"0000033e",x"00000340",
		x"00000342",x"00000344",x"00000346",x"00000348",x"0000034a",x"0000034c",x"0000034e",x"00000350",
		x"00000352",x"00000354",x"00000356",x"00000358",x"0000035a",x"0000035c",x"0000035e",x"00000360",
		x"00000362",x"00000364",x"00000366",x"00000368",x"0000036a",x"0000036c",x"0000036e",x"00000370",
		x"00000372",x"00000374",x"00000376",x"00000378",x"0000037a",x"0000037c",x"0000037e",x"00000380",
		x"00000382",x"00000384",x"00000386",x"00000388",x"0000038a",x"0000038c",x"0000038e",x"00000390",
		x"00000392",x"00000394",x"00000396",x"00000398",x"0000039a",x"0000039c",x"0000039e",x"000003a0",
		x"000003a2",x"000003a4",x"000003a6",x"000003a8",x"000003aa",x"000003ac",x"000003ae",x"000003b0",
		x"000003b2",x"000003b4",x"000003b6",x"000003b8",x"000003ba",x"000003bc",x"000003be",x"000003c0",
		x"000003c2",x"000003c4",x"000003c6",x"000003c8",x"000003ca",x"000003cc",x"000003ce",x"000003d0",
		x"000003d2",x"000003d4",x"000003d6",x"000003d8",x"000003da",x"000003dc",x"000003de",x"000003e0",
		x"000003e2",x"000003e4",x"000003e6",x"000003e8",x"000003ea",x"000003ec",x"000003ee",x"000003f0",
		x"000003f2",x"000003f4",x"000003f6",x"000003f8",x"000003fa",x"000003fc",x"000003fe",x"00000400",
		x"00000402",x"00000404",x"00000406",x"00000408",x"0000040a",x"0000040c",x"0000040e",x"00000410",
		x"00000412",x"00000414",x"00000416",x"00000418",x"0000041a",x"0000041c",x"0000041e",x"00000420",
		x"00000422",x"00000424",x"00000426",x"00000428",x"0000042a",x"0000042c",x"0000042e",x"00000430",
		x"00000432",x"00000434",x"00000436",x"00000438",x"0000043a",x"0000043c",x"0000043e",x"00000440",
		x"00000442",x"00000444",x"00000446",x"00000448",x"0000044a",x"0000044c",x"0000044e",x"00000450",
		x"00000452",x"00000454",x"00000456",x"00000458",x"0000045a",x"0000045c",x"0000045e",x"00000460",
		x"00000462",x"00000464",x"00000466",x"00000468",x"0000046a",x"0000046c",x"0000046e",x"00000470",
		x"00000472",x"00000474",x"00000476",x"00000478",x"0000047a",x"0000047c",x"0000047e",x"00000480",
		x"00000482",x"00000484",x"00000486",x"00000488",x"0000048a",x"0000048c",x"0000048e",x"00000490",
		x"00000492",x"00000494",x"00000496",x"00000498",x"0000049a",x"0000049c",x"0000049e",x"000004a0",
		x"000004a2",x"000004a4",x"000004a6",x"000004a8",x"000004aa",x"000004ac",x"000004ae",x"000004b0",
		x"000004b2",x"000004b4",x"000004b6",x"000004b8",x"000004ba",x"000004bc",x"000004be",x"000004c0",
		x"000004c2",x"000004c4",x"000004c6",x"000004c8",x"000004ca",x"000004cc",x"000004ce",x"000004d0",
		x"000004d2",x"000004d4",x"000004d6",x"000004d8",x"000004da",x"000004dc",x"000004de",x"000004e0",
		x"000004e2",x"000004e4",x"000004e6",x"000004e8",x"000004ea",x"000004ec",x"000004ee",x"000004f0",
		x"000004f2",x"000004f4",x"000004f6",x"000004f8",x"000004fa",x"000004fc",x"000004fe",x"00000500",
		x"00000502",x"00000504",x"00000506",x"00000508",x"0000050a",x"0000050c",x"0000050e",x"00000510",
		x"00000512",x"00000514",x"00000516",x"00000518",x"0000051a",x"0000051c",x"0000051e",x"00000520",
		x"00000522",x"00000524",x"00000526",x"00000528",x"0000052a",x"0000052c",x"0000052e",x"00000530",
		x"00000532",x"00000534",x"00000536",x"00000538",x"0000053a",x"0000053c",x"0000053e",x"00000540",
		x"00000542",x"00000544",x"00000546",x"00000548",x"0000054a",x"0000054c",x"0000054e",x"00000550",
		x"00000552",x"00000554",x"00000556",x"00000558",x"0000055a",x"0000055c",x"0000055e",x"00000560",
		x"00000562",x"00000564",x"00000566",x"00000568",x"0000056a",x"0000056c",x"0000056e",x"00000570",
		x"00000572",x"00000574",x"00000576",x"00000578",x"0000057a",x"0000057c",x"0000057e",x"00000580",
		x"00000582",x"00000584",x"00000586",x"00000588",x"0000058a",x"0000058c",x"0000058e",x"00000590",
		x"00000592",x"00000594",x"00000596",x"00000598",x"0000059a",x"0000059c",x"0000059e",x"000005a0",
		x"000005a2",x"000005a4",x"000005a6",x"000005a8",x"000005aa",x"000005ac",x"000005ae",x"000005b0",
		x"000005b2",x"000005b4",x"000005b6",x"000005b8",x"000005ba",x"000005bc",x"000005be",x"000005c0",
		x"000005c2",x"000005c4",x"000005c6",x"000005c8",x"000005ca",x"000005cc",x"000005ce",x"000005d0",
		x"000005d2",x"000005d4",x"000005d6",x"000005d8",x"000005da",x"000005dc",x"000005de",x"000005e0",
		x"000005e2",x"000005e4",x"000005e6",x"000005e8",x"000005ea",x"000005ec",x"000005ee",x"000005f0",
		x"000005f2",x"000005f4",x"000005f6",x"000005f8",x"000005fa",x"000005fc",x"000005fe",x"00000600",
		x"00000602",x"00000604",x"00000606",x"00000608",x"0000060a",x"0000060c",x"0000060e",x"00000610",
		x"00000612",x"00000614",x"00000616",x"00000618",x"0000061a",x"0000061c",x"0000061e",x"00000620",
		x"00000622",x"00000624",x"00000626",x"00000628",x"0000062a",x"0000062c",x"0000062e",x"00000630",
		x"00000632",x"00000634",x"00000636",x"00000638",x"0000063a",x"0000063c",x"0000063e",x"00000640",
		x"00000642",x"00000644",x"00000646",x"00000648",x"0000064a",x"0000064c",x"0000064e",x"00000650",
		x"00000652",x"00000654",x"00000656",x"00000658",x"0000065a",x"0000065c",x"0000065e",x"00000660",
		x"00000662",x"00000664",x"00000666",x"00000668",x"0000066a",x"0000066c",x"0000066e",x"00000670",
		x"00000672",x"00000674",x"00000676",x"00000678",x"0000067a",x"0000067c",x"0000067e",x"00000680",
		x"00000682",x"00000684",x"00000686",x"00000688",x"0000068a",x"0000068c",x"0000068e",x"00000690",
		x"00000692",x"00000694",x"00000696",x"00000698",x"0000069a",x"0000069c",x"0000069e",x"000006a0",
		x"000006a2",x"000006a4",x"000006a6",x"000006a8",x"000006aa",x"000006ac",x"000006ae",x"000006b0",
		x"000006b2",x"000006b4",x"000006b6",x"000006b8",x"000006ba",x"000006bc",x"000006be",x"000006c0",
		x"000006c2",x"000006c4",x"000006c6",x"000006c8",x"000006ca",x"000006cc",x"000006ce",x"000006d0",
		x"000006d2",x"000006d4",x"000006d6",x"000006d8",x"000006da",x"000006dc",x"000006de",x"000006e0",
		x"000006e2",x"000006e4",x"000006e6",x"000006e8",x"000006ea",x"000006ec",x"000006ee",x"000006f0",
		x"000006f2",x"000006f4",x"000006f6",x"000006f8",x"000006fa",x"000006fc",x"000006fe",x"00000700",
		x"00000702",x"00000704",x"00000706",x"00000708",x"0000070a",x"0000070c",x"0000070e",x"00000710",
		x"00000712",x"00000714",x"00000716",x"00000718",x"0000071a",x"0000071c",x"0000071e",x"00000720",
		x"00000722",x"00000724",x"00000726",x"00000728",x"0000072a",x"0000072c",x"0000072e",x"00000730",
		x"00000732",x"00000734",x"00000736",x"00000738",x"0000073a",x"0000073c",x"0000073e",x"00000740",
		x"00000742",x"00000744",x"00000746",x"00000748",x"0000074a",x"0000074c",x"0000074e",x"00000750",
		x"00000752",x"00000754",x"00000756",x"00000758",x"0000075a",x"0000075c",x"0000075e",x"00000760",
		x"00000762",x"00000764",x"00000766",x"00000768",x"0000076a",x"0000076c",x"0000076e",x"00000770",
		x"00000772",x"00000774",x"00000776",x"00000778",x"0000077a",x"0000077c",x"0000077e",x"00000780",
		x"00000782",x"00000784",x"00000786",x"00000788",x"0000078a",x"0000078c",x"0000078e",x"00000790",
		x"00000792",x"00000794",x"00000796",x"00000798",x"0000079a",x"0000079c",x"0000079e",x"000007a0",
		x"000007a2",x"000007a4",x"000007a6",x"000007a8",x"000007aa",x"000007ac",x"000007ae",x"000007b0",
		x"000007b2",x"000007b4",x"000007b6",x"000007b8",x"000007ba",x"000007bc",x"000007be",x"000007c0",
		x"000007c2",x"000007c4",x"000007c6",x"000007c8",x"000007ca",x"000007cc",x"000007ce",x"000007d0",
		x"000007d2",x"000007d4",x"000007d6",x"000007d8",x"000007da",x"000007dc",x"000007de",x"000007e0",
		x"000007e2",x"000007e4",x"000007e6",x"000007e8",x"000007ea",x"000007ec",x"000007ee",x"000007f0",
		x"000007f2",x"000007f4",x"000007f6",x"000007f8",x"000007fa",x"000007fc",x"000007fe",x"00000800",
		x"00000802",x"00000804",x"00000806",x"00000808",x"0000080a",x"0000080c",x"0000080e",x"00000810",
		x"00000812",x"00000814",x"00000816",x"00000818",x"0000081a",x"0000081c",x"0000081e",x"00000820",
		x"00000822",x"00000824",x"00000826",x"00000828",x"0000082a",x"0000082c",x"0000082e",x"00000830",
		x"00000832",x"00000834",x"00000836",x"00000838",x"0000083a",x"0000083c",x"0000083e",x"00000840",
		x"00000842",x"00000844",x"00000846",x"00000848",x"0000084a",x"0000084c",x"0000084e",x"00000850",
		x"00000852",x"00000854",x"00000856",x"00000858",x"0000085a",x"0000085c",x"0000085e",x"00000860",
		x"00000862",x"00000864",x"00000866",x"00000868",x"0000086a",x"0000086c",x"0000086e",x"00000870",
		x"00000872",x"00000874",x"00000876",x"00000878",x"0000087a",x"0000087c",x"0000087e",x"00000880",
		x"00000882",x"00000884",x"00000886",x"00000888",x"0000088a",x"0000088c",x"0000088e",x"00000890",
		x"00000892",x"00000894",x"00000896",x"00000898",x"0000089a",x"0000089c",x"0000089e",x"000008a0",
		x"000008a2",x"000008a4",x"000008a6",x"000008a8",x"000008aa",x"000008ac",x"000008ae",x"000008b0",
		x"000008b2",x"000008b4",x"000008b6",x"000008b8",x"000008ba",x"000008bc",x"000008be",x"000008c0",
		x"000008c2",x"000008c4",x"000008c6",x"000008c8",x"000008ca",x"000008cc",x"000008ce",x"000008d0",
		x"000008d2",x"000008d4",x"000008d6",x"000008d8",x"000008da",x"000008dc",x"000008de",x"000008e0",
		x"000008e2",x"000008e4",x"000008e6",x"000008e8",x"000008ea",x"000008ec",x"000008ee",x"000008f0",
		x"000008f2",x"000008f4",x"000008f6",x"000008f8",x"000008fa",x"000008fc",x"000008fe",x"00000900",
		x"00000902",x"00000904",x"00000906",x"00000908",x"0000090a",x"0000090c",x"0000090e",x"00000910",
		x"00000912",x"00000914",x"00000916",x"00000918",x"0000091a",x"0000091c",x"0000091e",x"00000920",
		x"00000922",x"00000924",x"00000926",x"00000928",x"0000092a",x"0000092c",x"0000092e",x"00000930",
		x"00000932",x"00000934",x"00000936",x"00000938",x"0000093a",x"0000093c",x"0000093e",x"00000940",
		x"00000942",x"00000944",x"00000946",x"00000948",x"0000094a",x"0000094c",x"0000094e",x"00000950",
		x"00000952",x"00000954",x"00000956",x"00000958",x"0000095a",x"0000095c",x"0000095e",x"00000960",
		x"00000962",x"00000964",x"00000966",x"00000968",x"0000096a",x"0000096c",x"0000096e",x"00000970",
		x"00000972",x"00000974",x"00000976",x"00000978",x"0000097a",x"0000097c",x"0000097e",x"00000980",
		x"00000982",x"00000984",x"00000986",x"00000988",x"0000098a",x"0000098c",x"0000098e",x"00000990",
		x"00000992",x"00000994",x"00000996",x"00000998",x"0000099a",x"0000099c",x"0000099e",x"000009a0",
		x"000009a2",x"000009a4",x"000009a6",x"000009a8",x"000009aa",x"000009ac",x"000009ae",x"000009b0",
		x"000009b2",x"000009b4",x"000009b6",x"000009b8",x"000009ba",x"000009bc",x"000009be",x"000009c0",
		x"000009c2",x"000009c4",x"000009c6",x"000009c8",x"000009ca",x"000009cc",x"000009ce",x"000009d0",
		x"000009d2",x"000009d4",x"000009d6",x"000009d8",x"000009da",x"000009dc",x"000009de",x"000009e0",
		x"000009e2",x"000009e4",x"000009e6",x"000009e8",x"000009ea",x"000009ec",x"000009ee",x"000009f0",
		x"000009f2",x"000009f4",x"000009f6",x"000009f8",x"000009fa",x"000009fc",x"000009fe",x"00000a00",
		x"00000a02",x"00000a04",x"00000a06",x"00000a08",x"00000a0a",x"00000a0c",x"00000a0e",x"00000a10",
		x"00000a12",x"00000a14",x"00000a16",x"00000a18",x"00000a1a",x"00000a1c",x"00000a1e",x"00000a20",
		x"00000a22",x"00000a24",x"00000a26",x"00000a28",x"00000a2a",x"00000a2c",x"00000a2e",x"00000a30",
		x"00000a32",x"00000a34",x"00000a36",x"00000a38",x"00000a3a",x"00000a3c",x"00000a3e",x"00000a40",
		x"00000a42",x"00000a44",x"00000a46",x"00000a48",x"00000a4a",x"00000a4c",x"00000a4e",x"00000a50",
		x"00000a52",x"00000a54",x"00000a56",x"00000a58",x"00000a5a",x"00000a5c",x"00000a5e",x"00000a60",
		x"00000a62",x"00000a64",x"00000a66",x"00000a68",x"00000a6a",x"00000a6c",x"00000a6e",x"00000a70",
		x"00000a72",x"00000a74",x"00000a76",x"00000a78",x"00000a7a",x"00000a7c",x"00000a7e",x"00000a80",
		x"00000a82",x"00000a84",x"00000a86",x"00000a88",x"00000a8a",x"00000a8c",x"00000a8e",x"00000a90",
		x"00000a92",x"00000a94",x"00000a96",x"00000a98",x"00000a9a",x"00000a9c",x"00000a9e",x"00000aa0",
		x"00000aa2",x"00000aa4",x"00000aa6",x"00000aa8",x"00000aaa",x"00000aac",x"00000aae",x"00000ab0",
		x"00000ab2",x"00000ab4",x"00000ab6",x"00000ab8",x"00000aba",x"00000abc",x"00000abe",x"00000ac0",
		x"00000ac2",x"00000ac4",x"00000ac6",x"00000ac8",x"00000aca",x"00000acc",x"00000ace",x"00000ad0",
		x"00000ad2",x"00000ad4",x"00000ad6",x"00000ad8",x"00000ada",x"00000adc",x"00000ade",x"00000ae0",
		x"00000ae2",x"00000ae4",x"00000ae6",x"00000ae8",x"00000aea",x"00000aec",x"00000aee",x"00000af0",
		x"00000af2",x"00000af4",x"00000af6",x"00000af8",x"00000afa",x"00000afc",x"00000afe",x"00000b00",
		x"00000b02",x"00000b04",x"00000b06",x"00000b08",x"00000b0a",x"00000b0c",x"00000b0e",x"00000b10",
		x"00000b12",x"00000b14",x"00000b16",x"00000b18",x"00000b1a",x"00000b1c",x"00000b1e",x"00000b20",
		x"00000b22",x"00000b24",x"00000b26",x"00000b28",x"00000b2a",x"00000b2c",x"00000b2e",x"00000b30",
		x"00000b32",x"00000b34",x"00000b36",x"00000b38",x"00000b3a",x"00000b3c",x"00000b3e",x"00000b40",
		x"00000b42",x"00000b44",x"00000b46",x"00000b48",x"00000b4a",x"00000b4c",x"00000b4e",x"00000b50",
		x"00000b52",x"00000b54",x"00000b56",x"00000b58",x"00000b5a",x"00000b5c",x"00000b5e",x"00000b60",
		x"00000b62",x"00000b64",x"00000b66",x"00000b68",x"00000b6a",x"00000b6c",x"00000b6e",x"00000b70",
		x"00000b72",x"00000b74",x"00000b76",x"00000b78",x"00000b7a",x"00000b7c",x"00000b7e",x"00000b80",
		x"00000b82",x"00000b84",x"00000b86",x"00000b88",x"00000b8a",x"00000b8c",x"00000b8e",x"00000b90",
		x"00000b92",x"00000b94",x"00000b96",x"00000b98",x"00000b9a",x"00000b9c",x"00000b9e",x"00000ba0",
		x"00000ba2",x"00000ba4",x"00000ba6",x"00000ba8",x"00000baa",x"00000bac",x"00000bae",x"00000bb0",
		x"00000bb2",x"00000bb4",x"00000bb6",x"00000bb8",x"00000bba",x"00000bbc",x"00000bbe",x"00000bc0",
		x"00000bc2",x"00000bc4",x"00000bc6",x"00000bc8",x"00000bca",x"00000bcc",x"00000bce",x"00000bd0",
		x"00000bd2",x"00000bd4",x"00000bd6",x"00000bd8",x"00000bda",x"00000bdc",x"00000bde",x"00000be0",
		x"00000be2",x"00000be4",x"00000be6",x"00000be8",x"00000bea",x"00000bec",x"00000bee",x"00000bf0",
		x"00000bf2",x"00000bf4",x"00000bf6",x"00000bf8",x"00000bfa",x"00000bfc",x"00000bfe",x"00000c00",
		x"00000c02",x"00000c04",x"00000c06",x"00000c08",x"00000c0a",x"00000c0c",x"00000c0e",x"00000c10",
		x"00000c12",x"00000c14",x"00000c16",x"00000c18",x"00000c1a",x"00000c1c",x"00000c1e",x"00000c20",
		x"00000c22",x"00000c24",x"00000c26",x"00000c28",x"00000c2a",x"00000c2c",x"00000c2e",x"00000c30",
		x"00000c32",x"00000c34",x"00000c36",x"00000c38",x"00000c3a",x"00000c3c",x"00000c3e",x"00000c40",
		x"00000c42",x"00000c44",x"00000c46",x"00000c48",x"00000c4a",x"00000c4c",x"00000c4e",x"00000c50",
		x"00000c52",x"00000c54",x"00000c56",x"00000c58",x"00000c5a",x"00000c5c",x"00000c5e",x"00000c60",
		x"00000c62",x"00000c64",x"00000c66",x"00000c68",x"00000c6a",x"00000c6c",x"00000c6e",x"00000c70",
		x"00000c72",x"00000c74",x"00000c76",x"00000c78",x"00000c7a",x"00000c7c",x"00000c7e",x"00000c80",
		x"00000c82",x"00000c84",x"00000c86",x"00000c88",x"00000c8a",x"00000c8c",x"00000c8e",x"00000c90",
		x"00000c92",x"00000c94",x"00000c96",x"00000c98",x"00000c9a",x"00000c9c",x"00000c9e",x"00000ca0",
		x"00000ca2",x"00000ca4",x"00000ca6",x"00000ca8",x"00000caa",x"00000cac",x"00000cae",x"00000cb0",
		x"00000cb2",x"00000cb4",x"00000cb6",x"00000cb8",x"00000cba",x"00000cbc",x"00000cbe",x"00000cc0",
		x"00000cc2",x"00000cc4",x"00000cc6",x"00000cc8",x"00000cca",x"00000ccc",x"00000cce",x"00000cd0",
		x"00000cd2",x"00000cd4",x"00000cd6",x"00000cd8",x"00000cda",x"00000cdc",x"00000cde",x"00000ce0",
		x"00000ce2",x"00000ce4",x"00000ce6",x"00000ce8",x"00000cea",x"00000cec",x"00000cee",x"00000cf0",
		x"00000cf2",x"00000cf4",x"00000cf6",x"00000cf8",x"00000cfa",x"00000cfc",x"00000cfe",x"00000d00",
		x"00000d02",x"00000d04",x"00000d06",x"00000d08",x"00000d0a",x"00000d0c",x"00000d0e",x"00000d10",
		x"00000d12",x"00000d14",x"00000d16",x"00000d18",x"00000d1a",x"00000d1c",x"00000d1e",x"00000d20",
		x"00000d22",x"00000d24",x"00000d26",x"00000d28",x"00000d2a",x"00000d2c",x"00000d2e",x"00000d30",
		x"00000d32",x"00000d34",x"00000d36",x"00000d38",x"00000d3a",x"00000d3c",x"00000d3e",x"00000d40",
		x"00000d42",x"00000d44",x"00000d46",x"00000d48",x"00000d4a",x"00000d4c",x"00000d4e",x"00000d50",
		x"00000d52",x"00000d54",x"00000d56",x"00000d58",x"00000d5a",x"00000d5c",x"00000d5e",x"00000d60",
		x"00000d62",x"00000d64",x"00000d66",x"00000d68",x"00000d6a",x"00000d6c",x"00000d6e",x"00000d70",
		x"00000d72",x"00000d74",x"00000d76",x"00000d78",x"00000d7a",x"00000d7c",x"00000d7e",x"00000d80",
		x"00000d82",x"00000d84",x"00000d86",x"00000d88",x"00000d8a",x"00000d8c",x"00000d8e",x"00000d90",
		x"00000d92",x"00000d94",x"00000d96",x"00000d98",x"00000d9a",x"00000d9c",x"00000d9e",x"00000da0",
		x"00000da2",x"00000da4",x"00000da6",x"00000da8",x"00000daa",x"00000dac",x"00000dae",x"00000db0",
		x"00000db2",x"00000db4",x"00000db6",x"00000db8",x"00000dba",x"00000dbc",x"00000dbe",x"00000dc0",
		x"00000dc2",x"00000dc4",x"00000dc6",x"00000dc8",x"00000dca",x"00000dcc",x"00000dce",x"00000dd0",
		x"00000dd2",x"00000dd4",x"00000dd6",x"00000dd8",x"00000dda",x"00000ddc",x"00000dde",x"00000de0",
		x"00000de2",x"00000de4",x"00000de6",x"00000de8",x"00000dea",x"00000dec",x"00000dee",x"00000df0",
		x"00000df2",x"00000df4",x"00000df6",x"00000df8",x"00000dfa",x"00000dfc",x"00000dfe",x"00000e00",
		x"00000e02",x"00000e04",x"00000e06",x"00000e08",x"00000e0a",x"00000e0c",x"00000e0e",x"00000e10",
		x"00000e12",x"00000e14",x"00000e16",x"00000e18",x"00000e1a",x"00000e1c",x"00000e1e",x"00000e20",
		x"00000e22",x"00000e24",x"00000e26",x"00000e28",x"00000e2a",x"00000e2c",x"00000e2e",x"00000e30",
		x"00000e32",x"00000e34",x"00000e36",x"00000e38",x"00000e3a",x"00000e3c",x"00000e3e",x"00000e40",
		x"00000e42",x"00000e44",x"00000e46",x"00000e48",x"00000e4a",x"00000e4c",x"00000e4e",x"00000e50",
		x"00000e52",x"00000e54",x"00000e56",x"00000e58",x"00000e5a",x"00000e5c",x"00000e5e",x"00000e60",
		x"00000e62",x"00000e64",x"00000e66",x"00000e68",x"00000e6a",x"00000e6c",x"00000e6e",x"00000e70",
		x"00000e72",x"00000e74",x"00000e76",x"00000e78",x"00000e7a",x"00000e7c",x"00000e7e",x"00000e80",
		x"00000e82",x"00000e84",x"00000e86",x"00000e88",x"00000e8a",x"00000e8c",x"00000e8e",x"00000e90",
		x"00000e92",x"00000e94",x"00000e96",x"00000e98",x"00000e9a",x"00000e9c",x"00000e9e",x"00000ea0",
		x"00000ea2",x"00000ea4",x"00000ea6",x"00000ea8",x"00000eaa",x"00000eac",x"00000eae",x"00000eb0",
		x"00000eb2",x"00000eb4",x"00000eb6",x"00000eb8",x"00000eba",x"00000ebc",x"00000ebe",x"00000ec0",
		x"00000ec2",x"00000ec4",x"00000ec6",x"00000ec8",x"00000eca",x"00000ecc",x"00000ece",x"00000ed0",
		x"00000ed2",x"00000ed4",x"00000ed6",x"00000ed8",x"00000eda",x"00000edc",x"00000ede",x"00000ee0",
		x"00000ee2",x"00000ee4",x"00000ee6",x"00000ee8",x"00000eea",x"00000eec",x"00000eee",x"00000ef0",
		x"00000ef2",x"00000ef4",x"00000ef6",x"00000ef8",x"00000efa",x"00000efc",x"00000efe",x"00000f00",
		x"00000f02",x"00000f04",x"00000f06",x"00000f08",x"00000f0a",x"00000f0c",x"00000f0e",x"00000f10",
		x"00000f12",x"00000f14",x"00000f16",x"00000f18",x"00000f1a",x"00000f1c",x"00000f1e",x"00000f20",
		x"00000f22",x"00000f24",x"00000f26",x"00000f28",x"00000f2a",x"00000f2c",x"00000f2e",x"00000f30",
		x"00000f32",x"00000f34",x"00000f36",x"00000f38",x"00000f3a",x"00000f3c",x"00000f3e",x"00000f40",
		x"00000f42",x"00000f44",x"00000f46",x"00000f48",x"00000f4a",x"00000f4c",x"00000f4e",x"00000f50",
		x"00000f52",x"00000f54",x"00000f56",x"00000f58",x"00000f5a",x"00000f5c",x"00000f5e",x"00000f60",
		x"00000f62",x"00000f64",x"00000f66",x"00000f68",x"00000f6a",x"00000f6c",x"00000f6e",x"00000f70",
		x"00000f72",x"00000f74",x"00000f76",x"00000f78",x"00000f7a",x"00000f7c",x"00000f7e",x"00000f80",
		x"00000f82",x"00000f84",x"00000f86",x"00000f88",x"00000f8a",x"00000f8c",x"00000f8e",x"00000f90",
		x"00000f92",x"00000f94",x"00000f96",x"00000f98",x"00000f9a",x"00000f9c",x"00000f9e",x"00000fa0",
		x"00000fa2",x"00000fa4",x"00000fa6",x"00000fa8",x"00000faa",x"00000fac",x"00000fae",x"00000fb0",
		x"00000fb2",x"00000fb4",x"00000fb6",x"00000fb8",x"00000fba",x"00000fbc",x"00000fbe",x"00000fc0",
		x"00000fc2",x"00000fc4",x"00000fc6",x"00000fc8",x"00000fca",x"00000fcc",x"00000fce",x"00000fd0",
		x"00000fd2",x"00000fd4",x"00000fd6",x"00000fd8",x"00000fda",x"00000fdc",x"00000fde",x"00000fe0",
		x"00000fe2",x"00000fe4",x"00000fe6",x"00000fe8",x"00000fea",x"00000fec",x"00000fee",x"00000ff0",
		x"00000ff2",x"00000ff4",x"00000ff6",x"00000ff8",x"00000ffa",x"00000ffc",x"00000ffe",x"00001000",
		x"00001002",x"00001004",x"00001006",x"00001008",x"0000100a",x"0000100c",x"0000100e",x"00001010",
		x"00001012",x"00001014",x"00001016",x"00001018",x"0000101a",x"0000101c",x"0000101e",x"00001020",
		x"00001022",x"00001024",x"00001026",x"00001028",x"0000102a",x"0000102c",x"0000102e",x"00001030",
		x"00001032",x"00001034",x"00001036",x"00001038",x"0000103a",x"0000103c",x"0000103e",x"00001040",
		x"00001042",x"00001044",x"00001046",x"00001048",x"0000104a",x"0000104c",x"0000104e",x"00001050",
		x"00001052",x"00001054",x"00001056",x"00001058",x"0000105a",x"0000105c",x"0000105e",x"00001060",
		x"00001062",x"00001064",x"00001066",x"00001068",x"0000106a",x"0000106c",x"0000106e",x"00001070",
		x"00001072",x"00001074",x"00001076",x"00001078",x"0000107a",x"0000107c",x"0000107e",x"00001080",
		x"00001082",x"00001084",x"00001086",x"00001088",x"0000108a",x"0000108c",x"0000108e",x"00001090",
		x"00001092",x"00001094",x"00001096",x"00001098",x"0000109a",x"0000109c",x"0000109e",x"000010a0",
		x"000010a2",x"000010a4",x"000010a6",x"000010a8",x"000010aa",x"000010ac",x"000010ae",x"000010b0",
		x"000010b2",x"000010b4",x"000010b6",x"000010b8",x"000010ba",x"000010bc",x"000010be",x"000010c0",
		x"000010c2",x"000010c4",x"000010c6",x"000010c8",x"000010ca",x"000010cc",x"000010ce",x"000010d0",
		x"000010d2",x"000010d4",x"000010d6",x"000010d8",x"000010da",x"000010dc",x"000010de",x"000010e0",
		x"000010e2",x"000010e4",x"000010e6",x"000010e8",x"000010ea",x"000010ec",x"000010ee",x"000010f0",
		x"000010f2",x"000010f4",x"000010f6",x"000010f8",x"000010fa",x"000010fc",x"000010fe",x"00001100",
		x"00001102",x"00001104",x"00001106",x"00001108",x"0000110a",x"0000110c",x"0000110e",x"00001110",
		x"00001112",x"00001114",x"00001116",x"00001118",x"0000111a",x"0000111c",x"0000111e",x"00001120",
		x"00001122",x"00001124",x"00001126",x"00001128",x"0000112a",x"0000112c",x"0000112e",x"00001130",
		x"00001132",x"00001134",x"00001136",x"00001138",x"0000113a",x"0000113c",x"0000113e",x"00001140",
		x"00001142",x"00001144",x"00001146",x"00001148",x"0000114a",x"0000114c",x"0000114e",x"00001150",
		x"00001152",x"00001154",x"00001156",x"00001158",x"0000115a",x"0000115c",x"0000115e",x"00001160",
		x"00001162",x"00001164",x"00001166",x"00001168",x"0000116a",x"0000116c",x"0000116e",x"00001170",
		x"00001172",x"00001174",x"00001176",x"00001178",x"0000117a",x"0000117c",x"0000117e",x"00001180",
		x"00001182",x"00001184",x"00001186",x"00001188",x"0000118a",x"0000118c",x"0000118e",x"00001190",
		x"00001192",x"00001194",x"00001196",x"00001198",x"0000119a",x"0000119c",x"0000119e",x"000011a0",
		x"000011a2",x"000011a4",x"000011a6",x"000011a8",x"000011aa",x"000011ac",x"000011ae",x"000011b0",
		x"000011b2",x"000011b4",x"000011b6",x"000011b8",x"000011ba",x"000011bc",x"000011be",x"000011c0",
		x"000011c2",x"000011c4",x"000011c6",x"000011c8",x"000011ca",x"000011cc",x"000011ce",x"000011d0",
		x"000011d2",x"000011d4",x"000011d6",x"000011d8",x"000011da",x"000011dc",x"000011de",x"000011e0",
		x"000011e2",x"000011e4",x"000011e6",x"000011e8",x"000011ea",x"000011ec",x"000011ee",x"000011f0",
		x"000011f2",x"000011f4",x"000011f6",x"000011f8",x"000011fa",x"000011fc",x"000011fe",x"00001200",
		x"00001202",x"00001204",x"00001206",x"00001208",x"0000120a",x"0000120c",x"0000120e",x"00001210",
		x"00001212",x"00001214",x"00001216",x"00001218",x"0000121a",x"0000121c",x"0000121e",x"00001220",
		x"00001222",x"00001224",x"00001226",x"00001228",x"0000122a",x"0000122c",x"0000122e",x"00001230",
		x"00001232",x"00001234",x"00001236",x"00001238",x"0000123a",x"0000123c",x"0000123e",x"00001240",
		x"00001242",x"00001244",x"00001246",x"00001248",x"0000124a",x"0000124c",x"0000124e",x"00001250",
		x"00001252",x"00001254",x"00001256",x"00001258",x"0000125a",x"0000125c",x"0000125e",x"00001260",
		x"00001262",x"00001264",x"00001266",x"00001268",x"0000126a",x"0000126c",x"0000126e",x"00001270",
		x"00001272",x"00001274",x"00001276",x"00001278",x"0000127a",x"0000127c",x"0000127e",x"00001280",
		x"00001282",x"00001284",x"00001286",x"00001288",x"0000128a",x"0000128c",x"0000128e",x"00001290",
		x"00001292",x"00001294",x"00001296",x"00001298",x"0000129a",x"0000129c",x"0000129e",x"000012a0",
		x"000012a2",x"000012a4",x"000012a6",x"000012a8",x"000012aa",x"000012ac",x"000012ae",x"000012b0",
		x"000012b2",x"000012b4",x"000012b6",x"000012b8",x"000012ba",x"000012bc",x"000012be",x"000012c0",
		x"000012c2",x"000012c4",x"000012c6",x"000012c8",x"000012ca",x"000012cc",x"000012ce",x"000012d0",
		x"000012d2",x"000012d4",x"000012d6",x"000012d8",x"000012da",x"000012dc",x"000012de",x"000012e0",
		x"000012e2",x"000012e4",x"000012e6",x"000012e8",x"000012ea",x"000012ec",x"000012ee",x"000012f0",
		x"000012f2",x"000012f4",x"000012f6",x"000012f8",x"000012fa",x"000012fc",x"000012fe",x"00001300",
		x"00001302",x"00001304",x"00001306",x"00001308",x"0000130a",x"0000130c",x"0000130e",x"00001310",
		x"00001312",x"00001314",x"00001316",x"00001318",x"0000131a",x"0000131c",x"0000131e",x"00001320",
		x"00001322",x"00001324",x"00001326",x"00001328",x"0000132a",x"0000132c",x"0000132e",x"00001330",
		x"00001332",x"00001334",x"00001336",x"00001338",x"0000133a",x"0000133c",x"0000133e",x"00001340",
		x"00001342",x"00001344",x"00001346",x"00001348",x"0000134a",x"0000134c",x"0000134e",x"00001350",
		x"00001352",x"00001354",x"00001356",x"00001358",x"0000135a",x"0000135c",x"0000135e",x"00001360",
		x"00001362",x"00001364",x"00001366",x"00001368",x"0000136a",x"0000136c",x"0000136e",x"00001370",
		x"00001372",x"00001374",x"00001376",x"00001378",x"0000137a",x"0000137c",x"0000137e",x"00001380",
		x"00001382",x"00001384",x"00001386",x"00001389",x"0000138b",x"0000138d",x"0000138f",x"00001391",
		x"00001393",x"00001395",x"00001397",x"00001399",x"0000139b",x"0000139d",x"0000139f",x"000013a1",
		x"000013a3",x"000013a5",x"000013a7",x"000013a9",x"000013ab",x"000013ad",x"000013af",x"000013b1",
		x"000013b3",x"000013b5",x"000013b7",x"000013b9",x"000013bb",x"000013bd",x"000013bf",x"000013c1",
		x"000013c3",x"000013c5",x"000013c7",x"000013c9",x"000013cb",x"000013cd",x"000013cf",x"000013d1",
		x"000013d3",x"000013d5",x"000013d7",x"000013d9",x"000013db",x"000013dd",x"000013df",x"000013e1",
		x"000013e3",x"000013e5",x"000013e7",x"000013e9",x"000013eb",x"000013ed",x"000013ef",x"000013f1",
		x"000013f3",x"000013f5",x"000013f7",x"000013f9",x"000013fb",x"000013fd",x"000013ff",x"00001401",
		x"00001403",x"00001405",x"00001407",x"00001409",x"0000140b",x"0000140d",x"0000140f",x"00001411",
		x"00001413",x"00001415",x"00001417",x"00001419",x"0000141b",x"0000141d",x"0000141f",x"00001421",
		x"00001423",x"00001425",x"00001427",x"00001429",x"0000142b",x"0000142d",x"0000142f",x"00001431",
		x"00001433",x"00001435",x"00001437",x"00001439",x"0000143b",x"0000143d",x"0000143f",x"00001441",
		x"00001443",x"00001445",x"00001447",x"00001449",x"0000144b",x"0000144d",x"0000144f",x"00001451",
		x"00001453",x"00001455",x"00001457",x"00001459",x"0000145b",x"0000145d",x"0000145f",x"00001461",
		x"00001463",x"00001465",x"00001467",x"00001469",x"0000146b",x"0000146d",x"0000146f",x"00001471",
		x"00001473",x"00001475",x"00001477",x"00001479",x"0000147b",x"0000147d",x"0000147f",x"00001481",
		x"00001483",x"00001485",x"00001487",x"00001489",x"0000148b",x"0000148d",x"0000148f",x"00001491",
		x"00001493",x"00001495",x"00001497",x"00001499",x"0000149b",x"0000149d",x"0000149f",x"000014a1",
		x"000014a3",x"000014a5",x"000014a7",x"000014a9",x"000014ab",x"000014ad",x"000014af",x"000014b1",
		x"000014b3",x"000014b5",x"000014b7",x"000014b9",x"000014bb",x"000014bd",x"000014bf",x"000014c1",
		x"000014c3",x"000014c5",x"000014c7",x"000014c9",x"000014cb",x"000014cd",x"000014cf",x"000014d1",
		x"000014d3",x"000014d5",x"000014d7",x"000014d9",x"000014db",x"000014dd",x"000014df",x"000014e1",
		x"000014e3",x"000014e5",x"000014e7",x"000014e9",x"000014eb",x"000014ed",x"000014ef",x"000014f1",
		x"000014f3",x"000014f5",x"000014f7",x"000014f9",x"000014fb",x"000014fd",x"000014ff",x"00001501",
		x"00001503",x"00001505",x"00001507",x"00001509",x"0000150b",x"0000150d",x"0000150f",x"00001511",
		x"00001513",x"00001515",x"00001517",x"00001519",x"0000151b",x"0000151d",x"0000151f",x"00001521",
		x"00001523",x"00001525",x"00001527",x"00001529",x"0000152b",x"0000152d",x"0000152f",x"00001531",
		x"00001533",x"00001535",x"00001537",x"00001539",x"0000153b",x"0000153d",x"0000153f",x"00001541",
		x"00001543",x"00001545",x"00001547",x"00001549",x"0000154b",x"0000154d",x"0000154f",x"00001551",
		x"00001553",x"00001555",x"00001557",x"00001559",x"0000155b",x"0000155d",x"0000155f",x"00001561",
		x"00001563",x"00001565",x"00001567",x"00001569",x"0000156b",x"0000156d",x"0000156f",x"00001571",
		x"00001573",x"00001575",x"00001577",x"00001579",x"0000157b",x"0000157d",x"0000157f",x"00001581",
		x"00001583",x"00001585",x"00001587",x"00001589",x"0000158b",x"0000158d",x"0000158f",x"00001591",
		x"00001593",x"00001595",x"00001597",x"00001599",x"0000159b",x"0000159d",x"0000159f",x"000015a1",
		x"000015a3",x"000015a5",x"000015a7",x"000015a9",x"000015ab",x"000015ad",x"000015af",x"000015b1",
		x"000015b3",x"000015b5",x"000015b7",x"000015b9",x"000015bb",x"000015bd",x"000015bf",x"000015c1",
		x"000015c3",x"000015c5",x"000015c7",x"000015c9",x"000015cb",x"000015cd",x"000015cf",x"000015d1",
		x"000015d3",x"000015d5",x"000015d7",x"000015d9",x"000015db",x"000015dd",x"000015df",x"000015e1",
		x"000015e3",x"000015e5",x"000015e7",x"000015e9",x"000015eb",x"000015ed",x"000015ef",x"000015f1",
		x"000015f3",x"000015f5",x"000015f7",x"000015f9",x"000015fb",x"000015fd",x"000015ff",x"00001601",
		x"00001603",x"00001605",x"00001607",x"00001609",x"0000160b",x"0000160d",x"0000160f",x"00001611",
		x"00001613",x"00001615",x"00001617",x"00001619",x"0000161b",x"0000161d",x"0000161f",x"00001621",
		x"00001623",x"00001625",x"00001627",x"00001629",x"0000162b",x"0000162d",x"0000162f",x"00001631",
		x"00001633",x"00001635",x"00001637",x"00001639",x"0000163b",x"0000163d",x"0000163f",x"00001641",
		x"00001643",x"00001645",x"00001647",x"00001649",x"0000164b",x"0000164d",x"0000164f",x"00001651",
		x"00001653",x"00001655",x"00001657",x"00001659",x"0000165b",x"0000165d",x"0000165f",x"00001661",
		x"00001663",x"00001665",x"00001667",x"00001669",x"0000166b",x"0000166d",x"0000166f",x"00001671",
		x"00001673",x"00001675",x"00001677",x"00001679",x"0000167b",x"0000167d",x"0000167f",x"00001681",
		x"00001683",x"00001685",x"00001687",x"00001689",x"0000168b",x"0000168d",x"0000168f",x"00001691",
		x"00001693",x"00001695",x"00001697",x"00001699",x"0000169b",x"0000169d",x"0000169f",x"000016a1",
		x"000016a3",x"000016a5",x"000016a7",x"000016a9",x"000016ab",x"000016ad",x"000016af",x"000016b1",
		x"000016b3",x"000016b5",x"000016b7",x"000016b9",x"000016bb",x"000016bd",x"000016bf",x"000016c1",
		x"000016c3",x"000016c5",x"000016c7",x"000016c9",x"000016cb",x"000016cd",x"000016cf",x"000016d1",
		x"000016d3",x"000016d5",x"000016d7",x"000016d9",x"000016db",x"000016dd",x"000016df",x"000016e1",
		x"000016e3",x"000016e5",x"000016e7",x"000016e9",x"000016eb",x"000016ed",x"000016ef",x"000016f1",
		x"000016f3",x"000016f5",x"000016f7",x"000016f9",x"000016fb",x"000016fd",x"000016ff",x"00001701",
		x"00001703",x"00001705",x"00001707",x"00001709",x"0000170b",x"0000170d",x"0000170f",x"00001711",
		x"00001713",x"00001715",x"00001717",x"00001719",x"0000171b",x"0000171d",x"0000171f",x"00001721",
		x"00001723",x"00001725",x"00001727",x"00001729",x"0000172b",x"0000172d",x"0000172f",x"00001731",
		x"00001733",x"00001735",x"00001737",x"00001739",x"0000173b",x"0000173d",x"0000173f",x"00001741",
		x"00001743",x"00001745",x"00001747",x"00001749",x"0000174b",x"0000174d",x"0000174f",x"00001751",
		x"00001753",x"00001755",x"00001757",x"00001759",x"0000175b",x"0000175d",x"0000175f",x"00001761",
		x"00001763",x"00001765",x"00001767",x"00001769",x"0000176b",x"0000176d",x"0000176f",x"00001771",
		x"00001773",x"00001775",x"00001777",x"00001779",x"0000177b",x"0000177d",x"0000177f",x"00001781",
		x"00001783",x"00001785",x"00001787",x"00001789",x"0000178b",x"0000178d",x"0000178f",x"00001791",
		x"00001793",x"00001795",x"00001797",x"00001799",x"0000179b",x"0000179d",x"0000179f",x"000017a1",
		x"000017a3",x"000017a5",x"000017a7",x"000017a9",x"000017ab",x"000017ad",x"000017af",x"000017b1",
		x"000017b3",x"000017b5",x"000017b7",x"000017b9",x"000017bb",x"000017bd",x"000017bf",x"000017c1",
		x"000017c3",x"000017c5",x"000017c7",x"000017c9",x"000017cb",x"000017cd",x"000017cf",x"000017d1",
		x"000017d3",x"000017d5",x"000017d7",x"000017d9",x"000017db",x"000017dd",x"000017df",x"000017e1",
		x"000017e3",x"000017e5",x"000017e7",x"000017e9",x"000017eb",x"000017ed",x"000017ef",x"000017f1",
		x"000017f3",x"000017f5",x"000017f7",x"000017f9",x"000017fb",x"000017fd",x"000017ff",x"00001801",
		x"00001803",x"00001805",x"00001807",x"00001809",x"0000180b",x"0000180d",x"0000180f",x"00001811",
		x"00001813",x"00001815",x"00001817",x"00001819",x"0000181b",x"0000181d",x"0000181f",x"00001821",
		x"00001823",x"00001825",x"00001827",x"00001829",x"0000182b",x"0000182d",x"0000182f",x"00001831",
		x"00001833",x"00001835",x"00001837",x"00001839",x"0000183b",x"0000183d",x"0000183f",x"00001841",
		x"00001843",x"00001845",x"00001847",x"00001849",x"0000184b",x"0000184d",x"0000184f",x"00001851",
		x"00001853",x"00001855",x"00001857",x"00001859",x"0000185b",x"0000185d",x"0000185f",x"00001861",
		x"00001863",x"00001865",x"00001867",x"00001869",x"0000186b",x"0000186d",x"0000186f",x"00001871",
		x"00001873",x"00001875",x"00001877",x"00001879",x"0000187b",x"0000187d",x"0000187f",x"00001881",
		x"00001883",x"00001885",x"00001887",x"00001889",x"0000188b",x"0000188d",x"0000188f",x"00001891",
		x"00001893",x"00001895",x"00001897",x"00001899",x"0000189b",x"0000189d",x"0000189f",x"000018a1",
		x"000018a3",x"000018a5",x"000018a7",x"000018a9",x"000018ab",x"000018ad",x"000018af",x"000018b1",
		x"000018b3",x"000018b5",x"000018b7",x"000018b9",x"000018bb",x"000018bd",x"000018bf",x"000018c1",
		x"000018c3",x"000018c5",x"000018c7",x"000018c9",x"000018cb",x"000018cd",x"000018cf",x"000018d1",
		x"000018d3",x"000018d5",x"000018d7",x"000018d9",x"000018db",x"000018dd",x"000018df",x"000018e1",
		x"000018e3",x"000018e5",x"000018e7",x"000018e9",x"000018eb",x"000018ed",x"000018ef",x"000018f1",
		x"000018f3",x"000018f5",x"000018f7",x"000018f9",x"000018fb",x"000018fd",x"000018ff",x"00001901",
		x"00001903",x"00001905",x"00001907",x"00001909",x"0000190b",x"0000190d",x"0000190f",x"00001911",
		x"00001913",x"00001915",x"00001917",x"00001919",x"0000191b",x"0000191d",x"0000191f",x"00001921",
		x"00001923",x"00001925",x"00001927",x"00001929",x"0000192b",x"0000192d",x"0000192f",x"00001931",
		x"00001933",x"00001935",x"00001937",x"00001939",x"0000193b",x"0000193d",x"0000193f",x"00001941",
		x"00001943",x"00001945",x"00001947",x"00001949",x"0000194b",x"0000194d",x"0000194f",x"00001951",
		x"00001953",x"00001955",x"00001957",x"00001959",x"0000195b",x"0000195d",x"0000195f",x"00001961",
		x"00001963",x"00001965",x"00001967",x"00001969",x"0000196b",x"0000196d",x"0000196f",x"00001971",
		x"00001973",x"00001975",x"00001977",x"00001979",x"0000197b",x"0000197d",x"0000197f",x"00001981",
		x"00001983",x"00001985",x"00001987",x"00001989",x"0000198b",x"0000198d",x"0000198f",x"00001991",
		x"00001993",x"00001995",x"00001997",x"00001999",x"0000199b",x"0000199d",x"0000199f",x"000019a1",
		x"000019a3",x"000019a5",x"000019a7",x"000019a9",x"000019ab",x"000019ad",x"000019af",x"000019b1",
		x"000019b3",x"000019b5",x"000019b7",x"000019b9",x"000019bb",x"000019bd",x"000019bf",x"000019c1",
		x"000019c3",x"000019c5",x"000019c7",x"000019c9",x"000019cb",x"000019cd",x"000019cf",x"000019d1",
		x"000019d3",x"000019d5",x"000019d7",x"000019d9",x"000019db",x"000019dd",x"000019df",x"000019e1",
		x"000019e3",x"000019e5",x"000019e7",x"000019e9",x"000019eb",x"000019ed",x"000019ef",x"000019f1",
		x"000019f3",x"000019f5",x"000019f7",x"000019f9",x"000019fb",x"000019fd",x"000019ff",x"00001a01",
		x"00001a03",x"00001a05",x"00001a07",x"00001a09",x"00001a0b",x"00001a0d",x"00001a0f",x"00001a11",
		x"00001a13",x"00001a15",x"00001a17",x"00001a19",x"00001a1b",x"00001a1d",x"00001a1f",x"00001a21",
		x"00001a23",x"00001a25",x"00001a27",x"00001a29",x"00001a2b",x"00001a2d",x"00001a2f",x"00001a31",
		x"00001a33",x"00001a35",x"00001a37",x"00001a39",x"00001a3b",x"00001a3d",x"00001a3f",x"00001a41",
		x"00001a43",x"00001a45",x"00001a47",x"00001a49",x"00001a4b",x"00001a4d",x"00001a4f",x"00001a51",
		x"00001a53",x"00001a55",x"00001a57",x"00001a59",x"00001a5b",x"00001a5d",x"00001a5f",x"00001a61",
		x"00001a63",x"00001a65",x"00001a67",x"00001a69",x"00001a6b",x"00001a6d",x"00001a6f",x"00001a71",
		x"00001a73",x"00001a75",x"00001a77",x"00001a79",x"00001a7b",x"00001a7d",x"00001a7f",x"00001a81",
		x"00001a83",x"00001a85",x"00001a87",x"00001a89",x"00001a8b",x"00001a8d",x"00001a8f",x"00001a91",
		x"00001a93",x"00001a95",x"00001a97",x"00001a99",x"00001a9b",x"00001a9d",x"00001a9f",x"00001aa1",
		x"00001aa3",x"00001aa5",x"00001aa7",x"00001aa9",x"00001aab",x"00001aad",x"00001aaf",x"00001ab1",
		x"00001ab3",x"00001ab5",x"00001ab7",x"00001ab9",x"00001abb",x"00001abd",x"00001abf",x"00001ac1",
		x"00001ac3",x"00001ac5",x"00001ac7",x"00001ac9",x"00001acb",x"00001acd",x"00001acf",x"00001ad1",
		x"00001ad3",x"00001ad5",x"00001ad7",x"00001ad9",x"00001adb",x"00001add",x"00001adf",x"00001ae1",
		x"00001ae3",x"00001ae5",x"00001ae7",x"00001ae9",x"00001aeb",x"00001aed",x"00001aef",x"00001af1",
		x"00001af3",x"00001af5",x"00001af7",x"00001af9",x"00001afb",x"00001afd",x"00001aff",x"00001b01",
		x"00001b03",x"00001b05",x"00001b07",x"00001b09",x"00001b0b",x"00001b0d",x"00001b0f",x"00001b11",
		x"00001b13",x"00001b15",x"00001b17",x"00001b19",x"00001b1b",x"00001b1d",x"00001b1f",x"00001b21",
		x"00001b23",x"00001b25",x"00001b27",x"00001b29",x"00001b2b",x"00001b2d",x"00001b2f",x"00001b31",
		x"00001b33",x"00001b35",x"00001b37",x"00001b39",x"00001b3b",x"00001b3d",x"00001b3f",x"00001b41",
		x"00001b43",x"00001b45",x"00001b47",x"00001b49",x"00001b4b",x"00001b4d",x"00001b4f",x"00001b51",
		x"00001b53",x"00001b55",x"00001b57",x"00001b59",x"00001b5b",x"00001b5d",x"00001b5f",x"00001b61",
		x"00001b63",x"00001b65",x"00001b67",x"00001b69",x"00001b6b",x"00001b6d",x"00001b6f",x"00001b71",
		x"00001b73",x"00001b75",x"00001b77",x"00001b79",x"00001b7b",x"00001b7d",x"00001b7f",x"00001b81",
		x"00001b83",x"00001b85",x"00001b87",x"00001b89",x"00001b8b",x"00001b8d",x"00001b8f",x"00001b91",
		x"00001b93",x"00001b95",x"00001b97",x"00001b99",x"00001b9b",x"00001b9d",x"00001b9f",x"00001ba1",
		x"00001ba3",x"00001ba5",x"00001ba7",x"00001ba9",x"00001bab",x"00001bad",x"00001baf",x"00001bb1",
		x"00001bb3",x"00001bb5",x"00001bb7",x"00001bb9",x"00001bbb",x"00001bbd",x"00001bbf",x"00001bc1",
		x"00001bc3",x"00001bc5",x"00001bc7",x"00001bc9",x"00001bcb",x"00001bcd",x"00001bcf",x"00001bd1",
		x"00001bd3",x"00001bd5",x"00001bd7",x"00001bd9",x"00001bdb",x"00001bdd",x"00001bdf",x"00001be1",
		x"00001be3",x"00001be5",x"00001be7",x"00001be9",x"00001beb",x"00001bed",x"00001bef",x"00001bf1",
		x"00001bf3",x"00001bf5",x"00001bf7",x"00001bf9",x"00001bfb",x"00001bfd",x"00001bff",x"00001c01",
		x"00001c03",x"00001c05",x"00001c07",x"00001c09",x"00001c0b",x"00001c0d",x"00001c0f",x"00001c11",
		x"00001c13",x"00001c15",x"00001c17",x"00001c19",x"00001c1b",x"00001c1d",x"00001c1f",x"00001c21",
		x"00001c23",x"00001c25",x"00001c27",x"00001c29",x"00001c2b",x"00001c2d",x"00001c2f",x"00001c31",
		x"00001c33",x"00001c35",x"00001c37",x"00001c39",x"00001c3b",x"00001c3d",x"00001c3f",x"00001c41",
		x"00001c43",x"00001c45",x"00001c47",x"00001c49",x"00001c4b",x"00001c4d",x"00001c4f",x"00001c51",
		x"00001c53",x"00001c55",x"00001c57",x"00001c59",x"00001c5b",x"00001c5d",x"00001c5f",x"00001c61",
		x"00001c63",x"00001c65",x"00001c67",x"00001c69",x"00001c6b",x"00001c6d",x"00001c6f",x"00001c71",
		x"00001c73",x"00001c75",x"00001c77",x"00001c79",x"00001c7b",x"00001c7d",x"00001c7f",x"00001c81",
		x"00001c83",x"00001c85",x"00001c87",x"00001c89",x"00001c8b",x"00001c8d",x"00001c8f",x"00001c91",
		x"00001c93",x"00001c95",x"00001c97",x"00001c99",x"00001c9b",x"00001c9d",x"00001c9f",x"00001ca1",
		x"00001ca3",x"00001ca5",x"00001ca7",x"00001ca9",x"00001cab",x"00001cad",x"00001caf",x"00001cb1",
		x"00001cb3",x"00001cb5",x"00001cb7",x"00001cb9",x"00001cbb",x"00001cbd",x"00001cbf",x"00001cc1",
		x"00001cc3",x"00001cc5",x"00001cc7",x"00001cc9",x"00001ccb",x"00001ccd",x"00001ccf",x"00001cd1",
		x"00001cd3",x"00001cd5",x"00001cd7",x"00001cd9",x"00001cdb",x"00001cdd",x"00001cdf",x"00001ce1",
		x"00001ce3",x"00001ce5",x"00001ce7",x"00001ce9",x"00001ceb",x"00001ced",x"00001cef",x"00001cf1",
		x"00001cf3",x"00001cf5",x"00001cf7",x"00001cf9",x"00001cfb",x"00001cfd",x"00001cff",x"00001d01",
		x"00001d03",x"00001d05",x"00001d07",x"00001d09",x"00001d0b",x"00001d0d",x"00001d0f",x"00001d11",
		x"00001d13",x"00001d15",x"00001d17",x"00001d19",x"00001d1b",x"00001d1d",x"00001d1f",x"00001d21",
		x"00001d23",x"00001d25",x"00001d27",x"00001d29",x"00001d2b",x"00001d2d",x"00001d2f",x"00001d31",
		x"00001d33",x"00001d35",x"00001d37",x"00001d39",x"00001d3b",x"00001d3d",x"00001d3f",x"00001d41",
		x"00001d43",x"00001d45",x"00001d47",x"00001d49",x"00001d4b",x"00001d4d",x"00001d4f",x"00001d51",
		x"00001d53",x"00001d55",x"00001d57",x"00001d59",x"00001d5b",x"00001d5d",x"00001d5f",x"00001d61",
		x"00001d63",x"00001d65",x"00001d67",x"00001d69",x"00001d6b",x"00001d6d",x"00001d6f",x"00001d71",
		x"00001d73",x"00001d75",x"00001d77",x"00001d79",x"00001d7b",x"00001d7d",x"00001d7f",x"00001d81",
		x"00001d83",x"00001d85",x"00001d87",x"00001d89",x"00001d8b",x"00001d8d",x"00001d8f",x"00001d91",
		x"00001d93",x"00001d95",x"00001d97",x"00001d99",x"00001d9b",x"00001d9d",x"00001d9f",x"00001da1",
		x"00001da3",x"00001da5",x"00001da7",x"00001da9",x"00001dab",x"00001dad",x"00001daf",x"00001db1",
		x"00001db3",x"00001db5",x"00001db7",x"00001db9",x"00001dbb",x"00001dbd",x"00001dbf",x"00001dc1",
		x"00001dc3",x"00001dc5",x"00001dc7",x"00001dc9",x"00001dcb",x"00001dcd",x"00001dcf",x"00001dd1",
		x"00001dd3",x"00001dd5",x"00001dd7",x"00001dd9",x"00001ddb",x"00001ddd",x"00001ddf",x"00001de1",
		x"00001de3",x"00001de5",x"00001de7",x"00001de9",x"00001deb",x"00001ded",x"00001def",x"00001df1",
		x"00001df3",x"00001df5",x"00001df7",x"00001df9",x"00001dfb",x"00001dfd",x"00001dff",x"00001e01",
		x"00001e03",x"00001e05",x"00001e07",x"00001e09",x"00001e0b",x"00001e0d",x"00001e0f",x"00001e11",
		x"00001e13",x"00001e15",x"00001e17",x"00001e19",x"00001e1b",x"00001e1d",x"00001e1f",x"00001e21",
		x"00001e23",x"00001e25",x"00001e27",x"00001e29",x"00001e2b",x"00001e2d",x"00001e2f",x"00001e31",
		x"00001e33",x"00001e35",x"00001e37",x"00001e39",x"00001e3b",x"00001e3d",x"00001e3f",x"00001e41",
		x"00001e43",x"00001e45",x"00001e47",x"00001e49",x"00001e4b",x"00001e4d",x"00001e4f",x"00001e51",
		x"00001e53",x"00001e55",x"00001e57",x"00001e59",x"00001e5b",x"00001e5d",x"00001e5f",x"00001e61",
		x"00001e63",x"00001e65",x"00001e67",x"00001e69",x"00001e6b",x"00001e6d",x"00001e6f",x"00001e71",
		x"00001e73",x"00001e75",x"00001e77",x"00001e79",x"00001e7b",x"00001e7d",x"00001e7f",x"00001e81",
		x"00001e83",x"00001e85",x"00001e87",x"00001e89",x"00001e8b",x"00001e8d",x"00001e8f",x"00001e91",
		x"00001e93",x"00001e95",x"00001e97",x"00001e99",x"00001e9b",x"00001e9d",x"00001e9f",x"00001ea1",
		x"00001ea3",x"00001ea5",x"00001ea7",x"00001ea9",x"00001eab",x"00001ead",x"00001eaf",x"00001eb1",
		x"00001eb3",x"00001eb5",x"00001eb7",x"00001eb9",x"00001ebb",x"00001ebd",x"00001ebf",x"00001ec1",
		x"00001ec3",x"00001ec5",x"00001ec7",x"00001ec9",x"00001ecb",x"00001ecd",x"00001ecf",x"00001ed1",
		x"00001ed3",x"00001ed5",x"00001ed7",x"00001ed9",x"00001edb",x"00001edd",x"00001edf",x"00001ee1",
		x"00001ee3",x"00001ee5",x"00001ee7",x"00001ee9",x"00001eeb",x"00001eed",x"00001eef",x"00001ef1",
		x"00001ef3",x"00001ef5",x"00001ef7",x"00001ef9",x"00001efb",x"00001efd",x"00001eff",x"00001f01",
		x"00001f03",x"00001f05",x"00001f07",x"00001f09",x"00001f0b",x"00001f0d",x"00001f0f",x"00001f11",
		x"00001f13",x"00001f15",x"00001f17",x"00001f19",x"00001f1b",x"00001f1d",x"00001f1f",x"00001f21",
		x"00001f23",x"00001f25",x"00001f27",x"00001f29",x"00001f2b",x"00001f2d",x"00001f2f",x"00001f31",
		x"00001f33",x"00001f35",x"00001f37",x"00001f39",x"00001f3b",x"00001f3d",x"00001f3f",x"00001f41",
		x"00001f43",x"00001f45",x"00001f47",x"00001f49",x"00001f4b",x"00001f4d",x"00001f4f",x"00001f51",
		x"00001f53",x"00001f55",x"00001f57",x"00001f59",x"00001f5b",x"00001f5d",x"00001f5f",x"00001f61",
		x"00001f63",x"00001f65",x"00001f67",x"00001f69",x"00001f6b",x"00001f6d",x"00001f6f",x"00001f71",
		x"00001f73",x"00001f75",x"00001f77",x"00001f79",x"00001f7b",x"00001f7d",x"00001f7f",x"00001f81",
		x"00001f83",x"00001f85",x"00001f87",x"00001f89",x"00001f8b",x"00001f8d",x"00001f8f",x"00001f91",
		x"00001f93",x"00001f95",x"00001f97",x"00001f99",x"00001f9b",x"00001f9d",x"00001f9f",x"00001fa1",
		x"00001fa3",x"00001fa5",x"00001fa7",x"00001fa9",x"00001fab",x"00001fad",x"00001faf",x"00001fb1",
		x"00001fb3",x"00001fb5",x"00001fb7",x"00001fb9",x"00001fbb",x"00001fbd",x"00001fbf",x"00001fc1",
		x"00001fc3",x"00001fc5",x"00001fc7",x"00001fc9",x"00001fcb",x"00001fcd",x"00001fcf",x"00001fd1",
		x"00001fd3",x"00001fd5",x"00001fd7",x"00001fd9",x"00001fdb",x"00001fdd",x"00001fdf",x"00001fe1",
		x"00001fe3",x"00001fe5",x"00001fe7",x"00001fe9",x"00001feb",x"00001fed",x"00001fef",x"00001ff1",
		x"00001ff3",x"00001ff5",x"00001ff7",x"00001ff9",x"00001ffb",x"00001ffd",x"00001fff",x"00002001",
		x"00002003",x"00002005",x"00002007",x"00002009",x"0000200b",x"0000200d",x"0000200f",x"00002011",
		x"00002013",x"00002015",x"00002017",x"00002019",x"0000201b",x"0000201d",x"0000201f",x"00002021",
		x"00002023",x"00002025",x"00002027",x"00002029",x"0000202b",x"0000202d",x"0000202f",x"00002031",
		x"00002033",x"00002035",x"00002037",x"00002039",x"0000203b",x"0000203d",x"0000203f",x"00002041",
		x"00002043",x"00002045",x"00002047",x"00002049",x"0000204b",x"0000204d",x"0000204f",x"00002051",
		x"00002053",x"00002055",x"00002057",x"00002059",x"0000205b",x"0000205d",x"0000205f",x"00002061",
		x"00002063",x"00002065",x"00002067",x"00002069",x"0000206b",x"0000206d",x"0000206f",x"00002071",
		x"00002073",x"00002075",x"00002077",x"00002079",x"0000207b",x"0000207d",x"0000207f",x"00002081",
		x"00002083",x"00002085",x"00002087",x"00002089",x"0000208b",x"0000208d",x"0000208f",x"00002091",
		x"00002093",x"00002095",x"00002097",x"00002099",x"0000209b",x"0000209d",x"0000209f",x"000020a1",
		x"000020a3",x"000020a5",x"000020a7",x"000020a9",x"000020ab",x"000020ad",x"000020af",x"000020b1",
		x"000020b3",x"000020b5",x"000020b7",x"000020b9",x"000020bb",x"000020bd",x"000020bf",x"000020c1",
		x"000020c3",x"000020c5",x"000020c7",x"000020c9",x"000020cb",x"000020cd",x"000020cf",x"000020d1",
		x"000020d3",x"000020d5",x"000020d7",x"000020d9",x"000020db",x"000020dd",x"000020df",x"000020e1",
		x"000020e3",x"000020e5",x"000020e7",x"000020e9",x"000020eb",x"000020ed",x"000020ef",x"000020f1",
		x"000020f3",x"000020f5",x"000020f7",x"000020f9",x"000020fb",x"000020fd",x"000020ff",x"00002101",
		x"00002103",x"00002105",x"00002107",x"00002109",x"0000210b",x"0000210d",x"0000210f",x"00002111",
		x"00002113",x"00002115",x"00002117",x"00002119",x"0000211b",x"0000211d",x"0000211f",x"00002121",
		x"00002123",x"00002125",x"00002127",x"00002129",x"0000212b",x"0000212d",x"0000212f",x"00002131",
		x"00002133",x"00002135",x"00002137",x"00002139",x"0000213b",x"0000213d",x"0000213f",x"00002141",
		x"00002143",x"00002145",x"00002147",x"00002149",x"0000214b",x"0000214d",x"0000214f",x"00002151",
		x"00002153",x"00002155",x"00002157",x"00002159",x"0000215b",x"0000215d",x"0000215f",x"00002161",
		x"00002163",x"00002165",x"00002167",x"00002169",x"0000216b",x"0000216d",x"0000216f",x"00002171",
		x"00002173",x"00002175",x"00002177",x"00002179",x"0000217b",x"0000217d",x"0000217f",x"00002181",
		x"00002183",x"00002185",x"00002187",x"00002189",x"0000218b",x"0000218d",x"0000218f",x"00002191",
		x"00002193",x"00002195",x"00002197",x"00002199",x"0000219b",x"0000219d",x"0000219f",x"000021a1",
		x"000021a3",x"000021a5",x"000021a7",x"000021a9",x"000021ab",x"000021ad",x"000021af",x"000021b1",
		x"000021b3",x"000021b5",x"000021b7",x"000021b9",x"000021bb",x"000021bd",x"000021bf",x"000021c1",
		x"000021c3",x"000021c5",x"000021c7",x"000021c9",x"000021cb",x"000021cd",x"000021cf",x"000021d1",
		x"000021d3",x"000021d5",x"000021d7",x"000021d9",x"000021db",x"000021dd",x"000021df",x"000021e1",
		x"000021e3",x"000021e5",x"000021e7",x"000021e9",x"000021eb",x"000021ed",x"000021ef",x"000021f1",
		x"000021f3",x"000021f5",x"000021f7",x"000021f9",x"000021fb",x"000021fd",x"000021ff",x"00002201",
		x"00002203",x"00002205",x"00002207",x"00002209",x"0000220b",x"0000220d",x"0000220f",x"00002211",
		x"00002213",x"00002215",x"00002217",x"00002219",x"0000221b",x"0000221d",x"0000221f",x"00002221",
		x"00002223",x"00002225",x"00002227",x"00002229",x"0000222b",x"0000222d",x"0000222f",x"00002231",
		x"00002233",x"00002235",x"00002237",x"00002239",x"0000223b",x"0000223d",x"0000223f",x"00002241",
		x"00002243",x"00002245",x"00002247",x"00002249",x"0000224b",x"0000224d",x"0000224f",x"00002251",
		x"00002253",x"00002255",x"00002257",x"00002259",x"0000225b",x"0000225d",x"0000225f",x"00002261",
		x"00002263",x"00002265",x"00002267",x"00002269",x"0000226b",x"0000226d",x"0000226f",x"00002271",
		x"00002273",x"00002275",x"00002277",x"00002279",x"0000227b",x"0000227d",x"0000227f",x"00002281",
		x"00002283",x"00002285",x"00002287",x"00002289",x"0000228b",x"0000228d",x"0000228f",x"00002291",
		x"00002293",x"00002295",x"00002297",x"00002299",x"0000229b",x"0000229d",x"0000229f",x"000022a1",
		x"000022a3",x"000022a5",x"000022a7",x"000022a9",x"000022ab",x"000022ad",x"000022af",x"000022b1",
		x"000022b3",x"000022b5",x"000022b7",x"000022b9",x"000022bb",x"000022bd",x"000022bf",x"000022c1",
		x"000022c3",x"000022c5",x"000022c7",x"000022c9",x"000022cb",x"000022cd",x"000022cf",x"000022d1",
		x"000022d3",x"000022d5",x"000022d7",x"000022d9",x"000022db",x"000022dd",x"000022df",x"000022e1",
		x"000022e3",x"000022e5",x"000022e7",x"000022e9",x"000022eb",x"000022ed",x"000022ef",x"000022f1",
		x"000022f3",x"000022f5",x"000022f7",x"000022f9",x"000022fb",x"000022fd",x"000022ff",x"00002301",
		x"00002303",x"00002305",x"00002307",x"00002309",x"0000230b",x"0000230d",x"0000230f",x"00002311",
		x"00002313",x"00002315",x"00002317",x"00002319",x"0000231b",x"0000231d",x"0000231f",x"00002321",
		x"00002323",x"00002325",x"00002327",x"00002329",x"0000232b",x"0000232d",x"0000232f",x"00002331",
		x"00002333",x"00002335",x"00002337",x"00002339",x"0000233b",x"0000233d",x"0000233f",x"00002341",
		x"00002343",x"00002345",x"00002347",x"00002349",x"0000234b",x"0000234d",x"0000234f",x"00002351",
		x"00002353",x"00002355",x"00002357",x"00002359",x"0000235b",x"0000235d",x"0000235f",x"00002361",
		x"00002363",x"00002365",x"00002367",x"00002369",x"0000236b",x"0000236d",x"0000236f",x"00002371",
		x"00002373",x"00002375",x"00002377",x"00002379",x"0000237b",x"0000237d",x"0000237f",x"00002381",
		x"00002383",x"00002385",x"00002387",x"00002389",x"0000238b",x"0000238d",x"0000238f",x"00002391",
		x"00002393",x"00002395",x"00002397",x"00002399",x"0000239b",x"0000239d",x"0000239f",x"000023a1",
		x"000023a3",x"000023a5",x"000023a7",x"000023a9",x"000023ab",x"000023ad",x"000023af",x"000023b1",
		x"000023b3",x"000023b5",x"000023b7",x"000023b9",x"000023bb",x"000023bd",x"000023bf",x"000023c1",
		x"000023c3",x"000023c5",x"000023c7",x"000023c9",x"000023cb",x"000023cd",x"000023cf",x"000023d1",
		x"000023d3",x"000023d5",x"000023d7",x"000023d9",x"000023db",x"000023dd",x"000023df",x"000023e1",
		x"000023e3",x"000023e5",x"000023e7",x"000023e9",x"000023eb",x"000023ed",x"000023ef",x"000023f1",
		x"000023f3",x"000023f5",x"000023f7",x"000023f9",x"000023fb",x"000023fd",x"000023ff",x"00002401",
		x"00002403",x"00002405",x"00002407",x"00002409",x"0000240b",x"0000240d",x"0000240f",x"00002411",
		x"00002413",x"00002415",x"00002417",x"00002419",x"0000241b",x"0000241d",x"0000241f",x"00002421",
		x"00002423",x"00002425",x"00002427",x"00002429",x"0000242b",x"0000242d",x"0000242f",x"00002431",
		x"00002433",x"00002435",x"00002437",x"00002439",x"0000243b",x"0000243d",x"0000243f",x"00002441",
		x"00002443",x"00002445",x"00002447",x"00002449",x"0000244b",x"0000244d",x"0000244f",x"00002451",
		x"00002453",x"00002455",x"00002457",x"00002459",x"0000245b",x"0000245d",x"0000245f",x"00002461",
		x"00002463",x"00002465",x"00002467",x"00002469",x"0000246b",x"0000246d",x"0000246f",x"00002471",
		x"00002473",x"00002475",x"00002477",x"00002479",x"0000247b",x"0000247d",x"0000247f",x"00002481",
		x"00002483",x"00002485",x"00002487",x"00002489",x"0000248b",x"0000248d",x"0000248f",x"00002491",
		x"00002493",x"00002495",x"00002497",x"00002499",x"0000249b",x"0000249d",x"0000249f",x"000024a1",
		x"000024a3",x"000024a5",x"000024a7",x"000024a9",x"000024ab",x"000024ad",x"000024af",x"000024b1",
		x"000024b3",x"000024b5",x"000024b7",x"000024b9",x"000024bb",x"000024bd",x"000024bf",x"000024c1",
		x"000024c3",x"000024c5",x"000024c7",x"000024c9",x"000024cb",x"000024cd",x"000024cf",x"000024d1",
		x"000024d3",x"000024d5",x"000024d7",x"000024d9",x"000024db",x"000024dd",x"000024df",x"000024e1",
		x"000024e3",x"000024e5",x"000024e7",x"000024e9",x"000024eb",x"000024ed",x"000024ef",x"000024f1",
		x"000024f3",x"000024f5",x"000024f7",x"000024f9",x"000024fb",x"000024fd",x"000024ff",x"00002501",
		x"00002503",x"00002505",x"00002507",x"00002509",x"0000250b",x"0000250d",x"0000250f",x"00002511",
		x"00002513",x"00002515",x"00002517",x"00002519",x"0000251b",x"0000251d",x"0000251f",x"00002521",
		x"00002523",x"00002525",x"00002527",x"00002529",x"0000252b",x"0000252d",x"0000252f",x"00002531",
		x"00002533",x"00002535",x"00002537",x"00002539",x"0000253b",x"0000253d",x"0000253f",x"00002541",
		x"00002543",x"00002545",x"00002547",x"00002549",x"0000254b",x"0000254d",x"0000254f",x"00002551",
		x"00002553",x"00002555",x"00002557",x"00002559",x"0000255b",x"0000255d",x"0000255f",x"00002561",
		x"00002563",x"00002565",x"00002567",x"00002569",x"0000256b",x"0000256d",x"0000256f",x"00002571",
		x"00002573",x"00002575",x"00002577",x"00002579",x"0000257b",x"0000257d",x"0000257f",x"00002581",
		x"00002583",x"00002585",x"00002587",x"00002589",x"0000258b",x"0000258d",x"0000258f",x"00002591",
		x"00002593",x"00002595",x"00002597",x"00002599",x"0000259b",x"0000259d",x"0000259f",x"000025a1",
		x"000025a3",x"000025a5",x"000025a7",x"000025a9",x"000025ab",x"000025ad",x"000025af",x"000025b1",
		x"000025b3",x"000025b5",x"000025b7",x"000025b9",x"000025bb",x"000025bd",x"000025bf",x"000025c1",
		x"000025c3",x"000025c5",x"000025c7",x"000025c9",x"000025cb",x"000025cd",x"000025cf",x"000025d1",
		x"000025d3",x"000025d5",x"000025d7",x"000025d9",x"000025db",x"000025dd",x"000025df",x"000025e1",
		x"000025e3",x"000025e5",x"000025e7",x"000025e9",x"000025eb",x"000025ed",x"000025ef",x"000025f1",
		x"000025f3",x"000025f5",x"000025f7",x"000025f9",x"000025fb",x"000025fd",x"000025ff",x"00002601",
		x"00002603",x"00002605",x"00002607",x"00002609",x"0000260b",x"0000260d",x"0000260f",x"00002611",
		x"00002613",x"00002615",x"00002617",x"00002619",x"0000261b",x"0000261d",x"0000261f",x"00002621",
		x"00002623",x"00002625",x"00002627",x"00002629",x"0000262b",x"0000262d",x"0000262f",x"00002631",
		x"00002633",x"00002635",x"00002637",x"00002639",x"0000263b",x"0000263d",x"0000263f",x"00002641",
		x"00002643",x"00002645",x"00002647",x"00002649",x"0000264b",x"0000264d",x"0000264f",x"00002651",
		x"00002653",x"00002655",x"00002657",x"00002659",x"0000265b",x"0000265d",x"0000265f",x"00002661",
		x"00002663",x"00002665",x"00002667",x"00002669",x"0000266b",x"0000266d",x"0000266f",x"00002671",
		x"00002673",x"00002675",x"00002677",x"00002679",x"0000267b",x"0000267d",x"0000267f",x"00002681",
		x"00002683",x"00002685",x"00002687",x"00002689",x"0000268b",x"0000268d",x"0000268f",x"00002691",
		x"00002693",x"00002695",x"00002697",x"00002699",x"0000269b",x"0000269d",x"0000269f",x"000026a1",
		x"000026a3",x"000026a5",x"000026a7",x"000026a9",x"000026ab",x"000026ad",x"000026af",x"000026b1",
		x"000026b3",x"000026b5",x"000026b7",x"000026b9",x"000026bb",x"000026bd",x"000026bf",x"000026c1",
		x"000026c3",x"000026c5",x"000026c7",x"000026c9",x"000026cb",x"000026cd",x"000026cf",x"000026d1",
		x"000026d3",x"000026d5",x"000026d7",x"000026d9",x"000026db",x"000026dd",x"000026df",x"000026e1",
		x"000026e3",x"000026e5",x"000026e7",x"000026e9",x"000026eb",x"000026ed",x"000026ef",x"000026f1",
		x"000026f3",x"000026f5",x"000026f7",x"000026f9",x"000026fb",x"000026fd",x"000026ff",x"00002701",
		x"00002703",x"00002705",x"00002707",x"00002709",x"0000270b",x"0000270d",x"0000270f",x"00002710",
		x"0000270f",x"0000270d",x"0000270b",x"00002709",x"00002707",x"00002705",x"00002703",x"00002701",
		x"000026ff",x"000026fd",x"000026fb",x"000026f9",x"000026f7",x"000026f5",x"000026f3",x"000026f1",
		x"000026ef",x"000026ed",x"000026eb",x"000026e9",x"000026e7",x"000026e5",x"000026e3",x"000026e1",
		x"000026df",x"000026dd",x"000026db",x"000026d9",x"000026d7",x"000026d5",x"000026d3",x"000026d1",
		x"000026cf",x"000026cd",x"000026cb",x"000026c9",x"000026c7",x"000026c5",x"000026c3",x"000026c1",
		x"000026bf",x"000026bd",x"000026bb",x"000026b9",x"000026b7",x"000026b5",x"000026b3",x"000026b1",
		x"000026af",x"000026ad",x"000026ab",x"000026a9",x"000026a7",x"000026a5",x"000026a3",x"000026a1",
		x"0000269f",x"0000269d",x"0000269b",x"00002699",x"00002697",x"00002695",x"00002693",x"00002691",
		x"0000268f",x"0000268d",x"0000268b",x"00002689",x"00002687",x"00002685",x"00002683",x"00002681",
		x"0000267f",x"0000267d",x"0000267b",x"00002679",x"00002677",x"00002675",x"00002673",x"00002671",
		x"0000266f",x"0000266d",x"0000266b",x"00002669",x"00002667",x"00002665",x"00002663",x"00002661",
		x"0000265f",x"0000265d",x"0000265b",x"00002659",x"00002657",x"00002655",x"00002653",x"00002651",
		x"0000264f",x"0000264d",x"0000264b",x"00002649",x"00002647",x"00002645",x"00002643",x"00002641",
		x"0000263f",x"0000263d",x"0000263b",x"00002639",x"00002637",x"00002635",x"00002633",x"00002631",
		x"0000262f",x"0000262d",x"0000262b",x"00002629",x"00002627",x"00002625",x"00002623",x"00002621",
		x"0000261f",x"0000261d",x"0000261b",x"00002619",x"00002617",x"00002615",x"00002613",x"00002611",
		x"0000260f",x"0000260d",x"0000260b",x"00002609",x"00002607",x"00002605",x"00002603",x"00002601",
		x"000025ff",x"000025fd",x"000025fb",x"000025f9",x"000025f7",x"000025f5",x"000025f3",x"000025f1",
		x"000025ef",x"000025ed",x"000025eb",x"000025e9",x"000025e7",x"000025e5",x"000025e3",x"000025e1",
		x"000025df",x"000025dd",x"000025db",x"000025d9",x"000025d7",x"000025d5",x"000025d3",x"000025d1",
		x"000025cf",x"000025cd",x"000025cb",x"000025c9",x"000025c7",x"000025c5",x"000025c3",x"000025c1",
		x"000025bf",x"000025bd",x"000025bb",x"000025b9",x"000025b7",x"000025b5",x"000025b3",x"000025b1",
		x"000025af",x"000025ad",x"000025ab",x"000025a9",x"000025a7",x"000025a5",x"000025a3",x"000025a1",
		x"0000259f",x"0000259d",x"0000259b",x"00002599",x"00002597",x"00002595",x"00002593",x"00002591",
		x"0000258f",x"0000258d",x"0000258b",x"00002589",x"00002587",x"00002585",x"00002583",x"00002581",
		x"0000257f",x"0000257d",x"0000257b",x"00002579",x"00002577",x"00002575",x"00002573",x"00002571",
		x"0000256f",x"0000256d",x"0000256b",x"00002569",x"00002567",x"00002565",x"00002563",x"00002561",
		x"0000255f",x"0000255d",x"0000255b",x"00002559",x"00002557",x"00002555",x"00002553",x"00002551",
		x"0000254f",x"0000254d",x"0000254b",x"00002549",x"00002547",x"00002545",x"00002543",x"00002541",
		x"0000253f",x"0000253d",x"0000253b",x"00002539",x"00002537",x"00002535",x"00002533",x"00002531",
		x"0000252f",x"0000252d",x"0000252b",x"00002529",x"00002527",x"00002525",x"00002523",x"00002521",
		x"0000251f",x"0000251d",x"0000251b",x"00002519",x"00002517",x"00002515",x"00002513",x"00002511",
		x"0000250f",x"0000250d",x"0000250b",x"00002509",x"00002507",x"00002505",x"00002503",x"00002501",
		x"000024ff",x"000024fd",x"000024fb",x"000024f9",x"000024f7",x"000024f5",x"000024f3",x"000024f1",
		x"000024ef",x"000024ed",x"000024eb",x"000024e9",x"000024e7",x"000024e5",x"000024e3",x"000024e1",
		x"000024df",x"000024dd",x"000024db",x"000024d9",x"000024d7",x"000024d5",x"000024d3",x"000024d1",
		x"000024cf",x"000024cd",x"000024cb",x"000024c9",x"000024c7",x"000024c5",x"000024c3",x"000024c1",
		x"000024bf",x"000024bd",x"000024bb",x"000024b9",x"000024b7",x"000024b5",x"000024b3",x"000024b1",
		x"000024af",x"000024ad",x"000024ab",x"000024a9",x"000024a7",x"000024a5",x"000024a3",x"000024a1",
		x"0000249f",x"0000249d",x"0000249b",x"00002499",x"00002497",x"00002495",x"00002493",x"00002491",
		x"0000248f",x"0000248d",x"0000248b",x"00002489",x"00002487",x"00002485",x"00002483",x"00002481",
		x"0000247f",x"0000247d",x"0000247b",x"00002479",x"00002477",x"00002475",x"00002473",x"00002471",
		x"0000246f",x"0000246d",x"0000246b",x"00002469",x"00002467",x"00002465",x"00002463",x"00002461",
		x"0000245f",x"0000245d",x"0000245b",x"00002459",x"00002457",x"00002455",x"00002453",x"00002451",
		x"0000244f",x"0000244d",x"0000244b",x"00002449",x"00002447",x"00002445",x"00002443",x"00002441",
		x"0000243f",x"0000243d",x"0000243b",x"00002439",x"00002437",x"00002435",x"00002433",x"00002431",
		x"0000242f",x"0000242d",x"0000242b",x"00002429",x"00002427",x"00002425",x"00002423",x"00002421",
		x"0000241f",x"0000241d",x"0000241b",x"00002419",x"00002417",x"00002415",x"00002413",x"00002411",
		x"0000240f",x"0000240d",x"0000240b",x"00002409",x"00002407",x"00002405",x"00002403",x"00002401",
		x"000023ff",x"000023fd",x"000023fb",x"000023f9",x"000023f7",x"000023f5",x"000023f3",x"000023f1",
		x"000023ef",x"000023ed",x"000023eb",x"000023e9",x"000023e7",x"000023e5",x"000023e3",x"000023e1",
		x"000023df",x"000023dd",x"000023db",x"000023d9",x"000023d7",x"000023d5",x"000023d3",x"000023d1",
		x"000023cf",x"000023cd",x"000023cb",x"000023c9",x"000023c7",x"000023c5",x"000023c3",x"000023c1",
		x"000023bf",x"000023bd",x"000023bb",x"000023b9",x"000023b7",x"000023b5",x"000023b3",x"000023b1",
		x"000023af",x"000023ad",x"000023ab",x"000023a9",x"000023a7",x"000023a5",x"000023a3",x"000023a1",
		x"0000239f",x"0000239d",x"0000239b",x"00002399",x"00002397",x"00002395",x"00002393",x"00002391",
		x"0000238f",x"0000238d",x"0000238b",x"00002389",x"00002387",x"00002385",x"00002383",x"00002381",
		x"0000237f",x"0000237d",x"0000237b",x"00002379",x"00002377",x"00002375",x"00002373",x"00002371",
		x"0000236f",x"0000236d",x"0000236b",x"00002369",x"00002367",x"00002365",x"00002363",x"00002361",
		x"0000235f",x"0000235d",x"0000235b",x"00002359",x"00002357",x"00002355",x"00002353",x"00002351",
		x"0000234f",x"0000234d",x"0000234b",x"00002349",x"00002347",x"00002345",x"00002343",x"00002341",
		x"0000233f",x"0000233d",x"0000233b",x"00002339",x"00002337",x"00002335",x"00002333",x"00002331",
		x"0000232f",x"0000232d",x"0000232b",x"00002329",x"00002327",x"00002325",x"00002323",x"00002321",
		x"0000231f",x"0000231d",x"0000231b",x"00002319",x"00002317",x"00002315",x"00002313",x"00002311",
		x"0000230f",x"0000230d",x"0000230b",x"00002309",x"00002307",x"00002305",x"00002303",x"00002301",
		x"000022ff",x"000022fd",x"000022fb",x"000022f9",x"000022f7",x"000022f5",x"000022f3",x"000022f1",
		x"000022ef",x"000022ed",x"000022eb",x"000022e9",x"000022e7",x"000022e5",x"000022e3",x"000022e1",
		x"000022df",x"000022dd",x"000022db",x"000022d9",x"000022d7",x"000022d5",x"000022d3",x"000022d1",
		x"000022cf",x"000022cd",x"000022cb",x"000022c9",x"000022c7",x"000022c5",x"000022c3",x"000022c1",
		x"000022bf",x"000022bd",x"000022bb",x"000022b9",x"000022b7",x"000022b5",x"000022b3",x"000022b1",
		x"000022af",x"000022ad",x"000022ab",x"000022a9",x"000022a7",x"000022a5",x"000022a3",x"000022a1",
		x"0000229f",x"0000229d",x"0000229b",x"00002299",x"00002297",x"00002295",x"00002293",x"00002291",
		x"0000228f",x"0000228d",x"0000228b",x"00002289",x"00002287",x"00002285",x"00002283",x"00002281",
		x"0000227f",x"0000227d",x"0000227b",x"00002279",x"00002277",x"00002275",x"00002273",x"00002271",
		x"0000226f",x"0000226d",x"0000226b",x"00002269",x"00002267",x"00002265",x"00002263",x"00002261",
		x"0000225f",x"0000225d",x"0000225b",x"00002259",x"00002257",x"00002255",x"00002253",x"00002251",
		x"0000224f",x"0000224d",x"0000224b",x"00002249",x"00002247",x"00002245",x"00002243",x"00002241",
		x"0000223f",x"0000223d",x"0000223b",x"00002239",x"00002237",x"00002235",x"00002233",x"00002231",
		x"0000222f",x"0000222d",x"0000222b",x"00002229",x"00002227",x"00002225",x"00002223",x"00002221",
		x"0000221f",x"0000221d",x"0000221b",x"00002219",x"00002217",x"00002215",x"00002213",x"00002211",
		x"0000220f",x"0000220d",x"0000220b",x"00002209",x"00002207",x"00002205",x"00002203",x"00002201",
		x"000021ff",x"000021fd",x"000021fb",x"000021f9",x"000021f7",x"000021f5",x"000021f3",x"000021f1",
		x"000021ef",x"000021ed",x"000021eb",x"000021e9",x"000021e7",x"000021e5",x"000021e3",x"000021e1",
		x"000021df",x"000021dd",x"000021db",x"000021d9",x"000021d7",x"000021d5",x"000021d3",x"000021d1",
		x"000021cf",x"000021cd",x"000021cb",x"000021c9",x"000021c7",x"000021c5",x"000021c3",x"000021c1",
		x"000021bf",x"000021bd",x"000021bb",x"000021b9",x"000021b7",x"000021b5",x"000021b3",x"000021b1",
		x"000021af",x"000021ad",x"000021ab",x"000021a9",x"000021a7",x"000021a5",x"000021a3",x"000021a1",
		x"0000219f",x"0000219d",x"0000219b",x"00002199",x"00002197",x"00002195",x"00002193",x"00002191",
		x"0000218f",x"0000218d",x"0000218b",x"00002189",x"00002187",x"00002185",x"00002183",x"00002181",
		x"0000217f",x"0000217d",x"0000217b",x"00002179",x"00002177",x"00002175",x"00002173",x"00002171",
		x"0000216f",x"0000216d",x"0000216b",x"00002169",x"00002167",x"00002165",x"00002163",x"00002161",
		x"0000215f",x"0000215d",x"0000215b",x"00002159",x"00002157",x"00002155",x"00002153",x"00002151",
		x"0000214f",x"0000214d",x"0000214b",x"00002149",x"00002147",x"00002145",x"00002143",x"00002141",
		x"0000213f",x"0000213d",x"0000213b",x"00002139",x"00002137",x"00002135",x"00002133",x"00002131",
		x"0000212f",x"0000212d",x"0000212b",x"00002129",x"00002127",x"00002125",x"00002123",x"00002121",
		x"0000211f",x"0000211d",x"0000211b",x"00002119",x"00002117",x"00002115",x"00002113",x"00002111",
		x"0000210f",x"0000210d",x"0000210b",x"00002109",x"00002107",x"00002105",x"00002103",x"00002101",
		x"000020ff",x"000020fd",x"000020fb",x"000020f9",x"000020f7",x"000020f5",x"000020f3",x"000020f1",
		x"000020ef",x"000020ed",x"000020eb",x"000020e9",x"000020e7",x"000020e5",x"000020e3",x"000020e1",
		x"000020df",x"000020dd",x"000020db",x"000020d9",x"000020d7",x"000020d5",x"000020d3",x"000020d1",
		x"000020cf",x"000020cd",x"000020cb",x"000020c9",x"000020c7",x"000020c5",x"000020c3",x"000020c1",
		x"000020bf",x"000020bd",x"000020bb",x"000020b9",x"000020b7",x"000020b5",x"000020b3",x"000020b1",
		x"000020af",x"000020ad",x"000020ab",x"000020a9",x"000020a7",x"000020a5",x"000020a3",x"000020a1",
		x"0000209f",x"0000209d",x"0000209b",x"00002099",x"00002097",x"00002095",x"00002093",x"00002091",
		x"0000208f",x"0000208d",x"0000208b",x"00002089",x"00002087",x"00002085",x"00002083",x"00002081",
		x"0000207f",x"0000207d",x"0000207b",x"00002079",x"00002077",x"00002075",x"00002073",x"00002071",
		x"0000206f",x"0000206d",x"0000206b",x"00002069",x"00002067",x"00002065",x"00002063",x"00002061",
		x"0000205f",x"0000205d",x"0000205b",x"00002059",x"00002057",x"00002055",x"00002053",x"00002051",
		x"0000204f",x"0000204d",x"0000204b",x"00002049",x"00002047",x"00002045",x"00002043",x"00002041",
		x"0000203f",x"0000203d",x"0000203b",x"00002039",x"00002037",x"00002035",x"00002033",x"00002031",
		x"0000202f",x"0000202d",x"0000202b",x"00002029",x"00002027",x"00002025",x"00002023",x"00002021",
		x"0000201f",x"0000201d",x"0000201b",x"00002019",x"00002017",x"00002015",x"00002013",x"00002011",
		x"0000200f",x"0000200d",x"0000200b",x"00002009",x"00002007",x"00002005",x"00002003",x"00002001",
		x"00001fff",x"00001ffd",x"00001ffb",x"00001ff9",x"00001ff7",x"00001ff5",x"00001ff3",x"00001ff1",
		x"00001fef",x"00001fed",x"00001feb",x"00001fe9",x"00001fe7",x"00001fe5",x"00001fe3",x"00001fe1",
		x"00001fdf",x"00001fdd",x"00001fdb",x"00001fd9",x"00001fd7",x"00001fd5",x"00001fd3",x"00001fd1",
		x"00001fcf",x"00001fcd",x"00001fcb",x"00001fc9",x"00001fc7",x"00001fc5",x"00001fc3",x"00001fc1",
		x"00001fbf",x"00001fbd",x"00001fbb",x"00001fb9",x"00001fb7",x"00001fb5",x"00001fb3",x"00001fb1",
		x"00001faf",x"00001fad",x"00001fab",x"00001fa9",x"00001fa7",x"00001fa5",x"00001fa3",x"00001fa1",
		x"00001f9f",x"00001f9d",x"00001f9b",x"00001f99",x"00001f97",x"00001f95",x"00001f93",x"00001f91",
		x"00001f8f",x"00001f8d",x"00001f8b",x"00001f89",x"00001f87",x"00001f85",x"00001f83",x"00001f81",
		x"00001f7f",x"00001f7d",x"00001f7b",x"00001f79",x"00001f77",x"00001f75",x"00001f73",x"00001f71",
		x"00001f6f",x"00001f6d",x"00001f6b",x"00001f69",x"00001f67",x"00001f65",x"00001f63",x"00001f61",
		x"00001f5f",x"00001f5d",x"00001f5b",x"00001f59",x"00001f57",x"00001f55",x"00001f53",x"00001f51",
		x"00001f4f",x"00001f4d",x"00001f4b",x"00001f49",x"00001f47",x"00001f45",x"00001f43",x"00001f41",
		x"00001f3f",x"00001f3d",x"00001f3b",x"00001f39",x"00001f37",x"00001f35",x"00001f33",x"00001f31",
		x"00001f2f",x"00001f2d",x"00001f2b",x"00001f29",x"00001f27",x"00001f25",x"00001f23",x"00001f21",
		x"00001f1f",x"00001f1d",x"00001f1b",x"00001f19",x"00001f17",x"00001f15",x"00001f13",x"00001f11",
		x"00001f0f",x"00001f0d",x"00001f0b",x"00001f09",x"00001f07",x"00001f05",x"00001f03",x"00001f01",
		x"00001eff",x"00001efd",x"00001efb",x"00001ef9",x"00001ef7",x"00001ef5",x"00001ef3",x"00001ef1",
		x"00001eef",x"00001eed",x"00001eeb",x"00001ee9",x"00001ee7",x"00001ee5",x"00001ee3",x"00001ee1",
		x"00001edf",x"00001edd",x"00001edb",x"00001ed9",x"00001ed7",x"00001ed5",x"00001ed3",x"00001ed1",
		x"00001ecf",x"00001ecd",x"00001ecb",x"00001ec9",x"00001ec7",x"00001ec5",x"00001ec3",x"00001ec1",
		x"00001ebf",x"00001ebd",x"00001ebb",x"00001eb9",x"00001eb7",x"00001eb5",x"00001eb3",x"00001eb1",
		x"00001eaf",x"00001ead",x"00001eab",x"00001ea9",x"00001ea7",x"00001ea5",x"00001ea3",x"00001ea1",
		x"00001e9f",x"00001e9d",x"00001e9b",x"00001e99",x"00001e97",x"00001e95",x"00001e93",x"00001e91",
		x"00001e8f",x"00001e8d",x"00001e8b",x"00001e89",x"00001e87",x"00001e85",x"00001e83",x"00001e81",
		x"00001e7f",x"00001e7d",x"00001e7b",x"00001e79",x"00001e77",x"00001e75",x"00001e73",x"00001e71",
		x"00001e6f",x"00001e6d",x"00001e6b",x"00001e69",x"00001e67",x"00001e65",x"00001e63",x"00001e61",
		x"00001e5f",x"00001e5d",x"00001e5b",x"00001e59",x"00001e57",x"00001e55",x"00001e53",x"00001e51",
		x"00001e4f",x"00001e4d",x"00001e4b",x"00001e49",x"00001e47",x"00001e45",x"00001e43",x"00001e41",
		x"00001e3f",x"00001e3d",x"00001e3b",x"00001e39",x"00001e37",x"00001e35",x"00001e33",x"00001e31",
		x"00001e2f",x"00001e2d",x"00001e2b",x"00001e29",x"00001e27",x"00001e25",x"00001e23",x"00001e21",
		x"00001e1f",x"00001e1d",x"00001e1b",x"00001e19",x"00001e17",x"00001e15",x"00001e13",x"00001e11",
		x"00001e0f",x"00001e0d",x"00001e0b",x"00001e09",x"00001e07",x"00001e05",x"00001e03",x"00001e01",
		x"00001dff",x"00001dfd",x"00001dfb",x"00001df9",x"00001df7",x"00001df5",x"00001df3",x"00001df1",
		x"00001def",x"00001ded",x"00001deb",x"00001de9",x"00001de7",x"00001de5",x"00001de3",x"00001de1",
		x"00001ddf",x"00001ddd",x"00001ddb",x"00001dd9",x"00001dd7",x"00001dd5",x"00001dd3",x"00001dd1",
		x"00001dcf",x"00001dcd",x"00001dcb",x"00001dc9",x"00001dc7",x"00001dc5",x"00001dc3",x"00001dc1",
		x"00001dbf",x"00001dbd",x"00001dbb",x"00001db9",x"00001db7",x"00001db5",x"00001db3",x"00001db1",
		x"00001daf",x"00001dad",x"00001dab",x"00001da9",x"00001da7",x"00001da5",x"00001da3",x"00001da1",
		x"00001d9f",x"00001d9d",x"00001d9b",x"00001d99",x"00001d97",x"00001d95",x"00001d93",x"00001d91",
		x"00001d8f",x"00001d8d",x"00001d8b",x"00001d89",x"00001d87",x"00001d85",x"00001d83",x"00001d81",
		x"00001d7f",x"00001d7d",x"00001d7b",x"00001d79",x"00001d77",x"00001d75",x"00001d73",x"00001d71",
		x"00001d6f",x"00001d6d",x"00001d6b",x"00001d69",x"00001d67",x"00001d65",x"00001d63",x"00001d61",
		x"00001d5f",x"00001d5d",x"00001d5b",x"00001d59",x"00001d57",x"00001d55",x"00001d53",x"00001d51",
		x"00001d4f",x"00001d4d",x"00001d4b",x"00001d49",x"00001d47",x"00001d45",x"00001d43",x"00001d41",
		x"00001d3f",x"00001d3d",x"00001d3b",x"00001d39",x"00001d37",x"00001d35",x"00001d33",x"00001d31",
		x"00001d2f",x"00001d2d",x"00001d2b",x"00001d29",x"00001d27",x"00001d25",x"00001d23",x"00001d21",
		x"00001d1f",x"00001d1d",x"00001d1b",x"00001d19",x"00001d17",x"00001d15",x"00001d13",x"00001d11",
		x"00001d0f",x"00001d0d",x"00001d0b",x"00001d09",x"00001d07",x"00001d05",x"00001d03",x"00001d01",
		x"00001cff",x"00001cfd",x"00001cfb",x"00001cf9",x"00001cf7",x"00001cf5",x"00001cf3",x"00001cf1",
		x"00001cef",x"00001ced",x"00001ceb",x"00001ce9",x"00001ce7",x"00001ce5",x"00001ce3",x"00001ce1",
		x"00001cdf",x"00001cdd",x"00001cdb",x"00001cd9",x"00001cd7",x"00001cd5",x"00001cd3",x"00001cd1",
		x"00001ccf",x"00001ccd",x"00001ccb",x"00001cc9",x"00001cc7",x"00001cc5",x"00001cc3",x"00001cc1",
		x"00001cbf",x"00001cbd",x"00001cbb",x"00001cb9",x"00001cb7",x"00001cb5",x"00001cb3",x"00001cb1",
		x"00001caf",x"00001cad",x"00001cab",x"00001ca9",x"00001ca7",x"00001ca5",x"00001ca3",x"00001ca1",
		x"00001c9f",x"00001c9d",x"00001c9b",x"00001c99",x"00001c97",x"00001c95",x"00001c93",x"00001c91",
		x"00001c8f",x"00001c8d",x"00001c8b",x"00001c89",x"00001c87",x"00001c85",x"00001c83",x"00001c81",
		x"00001c7f",x"00001c7d",x"00001c7b",x"00001c79",x"00001c77",x"00001c75",x"00001c73",x"00001c71",
		x"00001c6f",x"00001c6d",x"00001c6b",x"00001c69",x"00001c67",x"00001c65",x"00001c63",x"00001c61",
		x"00001c5f",x"00001c5d",x"00001c5b",x"00001c59",x"00001c57",x"00001c55",x"00001c53",x"00001c51",
		x"00001c4f",x"00001c4d",x"00001c4b",x"00001c49",x"00001c47",x"00001c45",x"00001c43",x"00001c41",
		x"00001c3f",x"00001c3d",x"00001c3b",x"00001c39",x"00001c37",x"00001c35",x"00001c33",x"00001c31",
		x"00001c2f",x"00001c2d",x"00001c2b",x"00001c29",x"00001c27",x"00001c25",x"00001c23",x"00001c21",
		x"00001c1f",x"00001c1d",x"00001c1b",x"00001c19",x"00001c17",x"00001c15",x"00001c13",x"00001c11",
		x"00001c0f",x"00001c0d",x"00001c0b",x"00001c09",x"00001c07",x"00001c05",x"00001c03",x"00001c01",
		x"00001bff",x"00001bfd",x"00001bfb",x"00001bf9",x"00001bf7",x"00001bf5",x"00001bf3",x"00001bf1",
		x"00001bef",x"00001bed",x"00001beb",x"00001be9",x"00001be7",x"00001be5",x"00001be3",x"00001be1",
		x"00001bdf",x"00001bdd",x"00001bdb",x"00001bd9",x"00001bd7",x"00001bd5",x"00001bd3",x"00001bd1",
		x"00001bcf",x"00001bcd",x"00001bcb",x"00001bc9",x"00001bc7",x"00001bc5",x"00001bc3",x"00001bc1",
		x"00001bbf",x"00001bbd",x"00001bbb",x"00001bb9",x"00001bb7",x"00001bb5",x"00001bb3",x"00001bb1",
		x"00001baf",x"00001bad",x"00001bab",x"00001ba9",x"00001ba7",x"00001ba5",x"00001ba3",x"00001ba1",
		x"00001b9f",x"00001b9d",x"00001b9b",x"00001b99",x"00001b97",x"00001b95",x"00001b93",x"00001b91",
		x"00001b8f",x"00001b8d",x"00001b8b",x"00001b89",x"00001b87",x"00001b85",x"00001b83",x"00001b81",
		x"00001b7f",x"00001b7d",x"00001b7b",x"00001b79",x"00001b77",x"00001b75",x"00001b73",x"00001b71",
		x"00001b6f",x"00001b6d",x"00001b6b",x"00001b69",x"00001b67",x"00001b65",x"00001b63",x"00001b61",
		x"00001b5f",x"00001b5d",x"00001b5b",x"00001b59",x"00001b57",x"00001b55",x"00001b53",x"00001b51",
		x"00001b4f",x"00001b4d",x"00001b4b",x"00001b49",x"00001b47",x"00001b45",x"00001b43",x"00001b41",
		x"00001b3f",x"00001b3d",x"00001b3b",x"00001b39",x"00001b37",x"00001b35",x"00001b33",x"00001b31",
		x"00001b2f",x"00001b2d",x"00001b2b",x"00001b29",x"00001b27",x"00001b25",x"00001b23",x"00001b21",
		x"00001b1f",x"00001b1d",x"00001b1b",x"00001b19",x"00001b17",x"00001b15",x"00001b13",x"00001b11",
		x"00001b0f",x"00001b0d",x"00001b0b",x"00001b09",x"00001b07",x"00001b05",x"00001b03",x"00001b01",
		x"00001aff",x"00001afd",x"00001afb",x"00001af9",x"00001af7",x"00001af5",x"00001af3",x"00001af1",
		x"00001aef",x"00001aed",x"00001aeb",x"00001ae9",x"00001ae7",x"00001ae5",x"00001ae3",x"00001ae1",
		x"00001adf",x"00001add",x"00001adb",x"00001ad9",x"00001ad7",x"00001ad5",x"00001ad3",x"00001ad1",
		x"00001acf",x"00001acd",x"00001acb",x"00001ac9",x"00001ac7",x"00001ac5",x"00001ac3",x"00001ac1",
		x"00001abf",x"00001abd",x"00001abb",x"00001ab9",x"00001ab7",x"00001ab5",x"00001ab3",x"00001ab1",
		x"00001aaf",x"00001aad",x"00001aab",x"00001aa9",x"00001aa7",x"00001aa5",x"00001aa3",x"00001aa1",
		x"00001a9f",x"00001a9d",x"00001a9b",x"00001a99",x"00001a97",x"00001a95",x"00001a93",x"00001a91",
		x"00001a8f",x"00001a8d",x"00001a8b",x"00001a89",x"00001a87",x"00001a85",x"00001a83",x"00001a81",
		x"00001a7f",x"00001a7d",x"00001a7b",x"00001a79",x"00001a77",x"00001a75",x"00001a73",x"00001a71",
		x"00001a6f",x"00001a6d",x"00001a6b",x"00001a69",x"00001a67",x"00001a65",x"00001a63",x"00001a61",
		x"00001a5f",x"00001a5d",x"00001a5b",x"00001a59",x"00001a57",x"00001a55",x"00001a53",x"00001a51",
		x"00001a4f",x"00001a4d",x"00001a4b",x"00001a49",x"00001a47",x"00001a45",x"00001a43",x"00001a41",
		x"00001a3f",x"00001a3d",x"00001a3b",x"00001a39",x"00001a37",x"00001a35",x"00001a33",x"00001a31",
		x"00001a2f",x"00001a2d",x"00001a2b",x"00001a29",x"00001a27",x"00001a25",x"00001a23",x"00001a21",
		x"00001a1f",x"00001a1d",x"00001a1b",x"00001a19",x"00001a17",x"00001a15",x"00001a13",x"00001a11",
		x"00001a0f",x"00001a0d",x"00001a0b",x"00001a09",x"00001a07",x"00001a05",x"00001a03",x"00001a01",
		x"000019ff",x"000019fd",x"000019fb",x"000019f9",x"000019f7",x"000019f5",x"000019f3",x"000019f1",
		x"000019ef",x"000019ed",x"000019eb",x"000019e9",x"000019e7",x"000019e5",x"000019e3",x"000019e1",
		x"000019df",x"000019dd",x"000019db",x"000019d9",x"000019d7",x"000019d5",x"000019d3",x"000019d1",
		x"000019cf",x"000019cd",x"000019cb",x"000019c9",x"000019c7",x"000019c5",x"000019c3",x"000019c1",
		x"000019bf",x"000019bd",x"000019bb",x"000019b9",x"000019b7",x"000019b5",x"000019b3",x"000019b1",
		x"000019af",x"000019ad",x"000019ab",x"000019a9",x"000019a7",x"000019a5",x"000019a3",x"000019a1",
		x"0000199f",x"0000199d",x"0000199b",x"00001999",x"00001997",x"00001995",x"00001993",x"00001991",
		x"0000198f",x"0000198d",x"0000198b",x"00001989",x"00001987",x"00001985",x"00001983",x"00001981",
		x"0000197f",x"0000197d",x"0000197b",x"00001979",x"00001977",x"00001975",x"00001973",x"00001971",
		x"0000196f",x"0000196d",x"0000196b",x"00001969",x"00001967",x"00001965",x"00001963",x"00001961",
		x"0000195f",x"0000195d",x"0000195b",x"00001959",x"00001957",x"00001955",x"00001953",x"00001951",
		x"0000194f",x"0000194d",x"0000194b",x"00001949",x"00001947",x"00001945",x"00001943",x"00001941",
		x"0000193f",x"0000193d",x"0000193b",x"00001939",x"00001937",x"00001935",x"00001933",x"00001931",
		x"0000192f",x"0000192d",x"0000192b",x"00001929",x"00001927",x"00001925",x"00001923",x"00001921",
		x"0000191f",x"0000191d",x"0000191b",x"00001919",x"00001917",x"00001915",x"00001913",x"00001911",
		x"0000190f",x"0000190d",x"0000190b",x"00001909",x"00001907",x"00001905",x"00001903",x"00001901",
		x"000018ff",x"000018fd",x"000018fb",x"000018f9",x"000018f7",x"000018f5",x"000018f3",x"000018f1",
		x"000018ef",x"000018ed",x"000018eb",x"000018e9",x"000018e7",x"000018e5",x"000018e3",x"000018e1",
		x"000018df",x"000018dd",x"000018db",x"000018d9",x"000018d7",x"000018d5",x"000018d3",x"000018d1",
		x"000018cf",x"000018cd",x"000018cb",x"000018c9",x"000018c7",x"000018c5",x"000018c3",x"000018c1",
		x"000018bf",x"000018bd",x"000018bb",x"000018b9",x"000018b7",x"000018b5",x"000018b3",x"000018b1",
		x"000018af",x"000018ad",x"000018ab",x"000018a9",x"000018a7",x"000018a5",x"000018a3",x"000018a1",
		x"0000189f",x"0000189d",x"0000189b",x"00001899",x"00001897",x"00001895",x"00001893",x"00001891",
		x"0000188f",x"0000188d",x"0000188b",x"00001889",x"00001887",x"00001885",x"00001883",x"00001881",
		x"0000187f",x"0000187d",x"0000187b",x"00001879",x"00001877",x"00001875",x"00001873",x"00001871",
		x"0000186f",x"0000186d",x"0000186b",x"00001869",x"00001867",x"00001865",x"00001863",x"00001861",
		x"0000185f",x"0000185d",x"0000185b",x"00001859",x"00001857",x"00001855",x"00001853",x"00001851",
		x"0000184f",x"0000184d",x"0000184b",x"00001849",x"00001847",x"00001845",x"00001843",x"00001841",
		x"0000183f",x"0000183d",x"0000183b",x"00001839",x"00001837",x"00001835",x"00001833",x"00001831",
		x"0000182f",x"0000182d",x"0000182b",x"00001829",x"00001827",x"00001825",x"00001823",x"00001821",
		x"0000181f",x"0000181d",x"0000181b",x"00001819",x"00001817",x"00001815",x"00001813",x"00001811",
		x"0000180f",x"0000180d",x"0000180b",x"00001809",x"00001807",x"00001805",x"00001803",x"00001801",
		x"000017ff",x"000017fd",x"000017fb",x"000017f9",x"000017f7",x"000017f5",x"000017f3",x"000017f1",
		x"000017ef",x"000017ed",x"000017eb",x"000017e9",x"000017e7",x"000017e5",x"000017e3",x"000017e1",
		x"000017df",x"000017dd",x"000017db",x"000017d9",x"000017d7",x"000017d5",x"000017d3",x"000017d1",
		x"000017cf",x"000017cd",x"000017cb",x"000017c9",x"000017c7",x"000017c5",x"000017c3",x"000017c1",
		x"000017bf",x"000017bd",x"000017bb",x"000017b9",x"000017b7",x"000017b5",x"000017b3",x"000017b1",
		x"000017af",x"000017ad",x"000017ab",x"000017a9",x"000017a7",x"000017a5",x"000017a3",x"000017a1",
		x"0000179f",x"0000179d",x"0000179b",x"00001799",x"00001797",x"00001795",x"00001793",x"00001791",
		x"0000178f",x"0000178d",x"0000178b",x"00001789",x"00001787",x"00001785",x"00001783",x"00001781",
		x"0000177f",x"0000177d",x"0000177b",x"00001779",x"00001777",x"00001775",x"00001773",x"00001771",
		x"0000176f",x"0000176d",x"0000176b",x"00001769",x"00001767",x"00001765",x"00001763",x"00001761",
		x"0000175f",x"0000175d",x"0000175b",x"00001759",x"00001757",x"00001755",x"00001753",x"00001751",
		x"0000174f",x"0000174d",x"0000174b",x"00001749",x"00001747",x"00001745",x"00001743",x"00001741",
		x"0000173f",x"0000173d",x"0000173b",x"00001739",x"00001737",x"00001735",x"00001733",x"00001731",
		x"0000172f",x"0000172d",x"0000172b",x"00001729",x"00001727",x"00001725",x"00001723",x"00001721",
		x"0000171f",x"0000171d",x"0000171b",x"00001719",x"00001717",x"00001715",x"00001713",x"00001711",
		x"0000170f",x"0000170d",x"0000170b",x"00001709",x"00001707",x"00001705",x"00001703",x"00001701",
		x"000016ff",x"000016fd",x"000016fb",x"000016f9",x"000016f7",x"000016f5",x"000016f3",x"000016f1",
		x"000016ef",x"000016ed",x"000016eb",x"000016e9",x"000016e7",x"000016e5",x"000016e3",x"000016e1",
		x"000016df",x"000016dd",x"000016db",x"000016d9",x"000016d7",x"000016d5",x"000016d3",x"000016d1",
		x"000016cf",x"000016cd",x"000016cb",x"000016c9",x"000016c7",x"000016c5",x"000016c3",x"000016c1",
		x"000016bf",x"000016bd",x"000016bb",x"000016b9",x"000016b7",x"000016b5",x"000016b3",x"000016b1",
		x"000016af",x"000016ad",x"000016ab",x"000016a9",x"000016a7",x"000016a5",x"000016a3",x"000016a1",
		x"0000169f",x"0000169d",x"0000169b",x"00001699",x"00001697",x"00001695",x"00001693",x"00001691",
		x"0000168f",x"0000168d",x"0000168b",x"00001689",x"00001687",x"00001685",x"00001683",x"00001681",
		x"0000167f",x"0000167d",x"0000167b",x"00001679",x"00001677",x"00001675",x"00001673",x"00001671",
		x"0000166f",x"0000166d",x"0000166b",x"00001669",x"00001667",x"00001665",x"00001663",x"00001661",
		x"0000165f",x"0000165d",x"0000165b",x"00001659",x"00001657",x"00001655",x"00001653",x"00001651",
		x"0000164f",x"0000164d",x"0000164b",x"00001649",x"00001647",x"00001645",x"00001643",x"00001641",
		x"0000163f",x"0000163d",x"0000163b",x"00001639",x"00001637",x"00001635",x"00001633",x"00001631",
		x"0000162f",x"0000162d",x"0000162b",x"00001629",x"00001627",x"00001625",x"00001623",x"00001621",
		x"0000161f",x"0000161d",x"0000161b",x"00001619",x"00001617",x"00001615",x"00001613",x"00001611",
		x"0000160f",x"0000160d",x"0000160b",x"00001609",x"00001607",x"00001605",x"00001603",x"00001601",
		x"000015ff",x"000015fd",x"000015fb",x"000015f9",x"000015f7",x"000015f5",x"000015f3",x"000015f1",
		x"000015ef",x"000015ed",x"000015eb",x"000015e9",x"000015e7",x"000015e5",x"000015e3",x"000015e1",
		x"000015df",x"000015dd",x"000015db",x"000015d9",x"000015d7",x"000015d5",x"000015d3",x"000015d1",
		x"000015cf",x"000015cd",x"000015cb",x"000015c9",x"000015c7",x"000015c5",x"000015c3",x"000015c1",
		x"000015bf",x"000015bd",x"000015bb",x"000015b9",x"000015b7",x"000015b5",x"000015b3",x"000015b1",
		x"000015af",x"000015ad",x"000015ab",x"000015a9",x"000015a7",x"000015a5",x"000015a3",x"000015a1",
		x"0000159f",x"0000159d",x"0000159b",x"00001599",x"00001597",x"00001595",x"00001593",x"00001591",
		x"0000158f",x"0000158d",x"0000158b",x"00001589",x"00001587",x"00001585",x"00001583",x"00001581",
		x"0000157f",x"0000157d",x"0000157b",x"00001579",x"00001577",x"00001575",x"00001573",x"00001571",
		x"0000156f",x"0000156d",x"0000156b",x"00001569",x"00001567",x"00001565",x"00001563",x"00001561",
		x"0000155f",x"0000155d",x"0000155b",x"00001559",x"00001557",x"00001555",x"00001553",x"00001551",
		x"0000154f",x"0000154d",x"0000154b",x"00001549",x"00001547",x"00001545",x"00001543",x"00001541",
		x"0000153f",x"0000153d",x"0000153b",x"00001539",x"00001537",x"00001535",x"00001533",x"00001531",
		x"0000152f",x"0000152d",x"0000152b",x"00001529",x"00001527",x"00001525",x"00001523",x"00001521",
		x"0000151f",x"0000151d",x"0000151b",x"00001519",x"00001517",x"00001515",x"00001513",x"00001511",
		x"0000150f",x"0000150d",x"0000150b",x"00001509",x"00001507",x"00001505",x"00001503",x"00001501",
		x"000014ff",x"000014fd",x"000014fb",x"000014f9",x"000014f7",x"000014f5",x"000014f3",x"000014f1",
		x"000014ef",x"000014ed",x"000014eb",x"000014e9",x"000014e7",x"000014e5",x"000014e3",x"000014e1",
		x"000014df",x"000014dd",x"000014db",x"000014d9",x"000014d7",x"000014d5",x"000014d3",x"000014d1",
		x"000014cf",x"000014cd",x"000014cb",x"000014c9",x"000014c7",x"000014c5",x"000014c3",x"000014c1",
		x"000014bf",x"000014bd",x"000014bb",x"000014b9",x"000014b7",x"000014b5",x"000014b3",x"000014b1",
		x"000014af",x"000014ad",x"000014ab",x"000014a9",x"000014a7",x"000014a5",x"000014a3",x"000014a1",
		x"0000149f",x"0000149d",x"0000149b",x"00001499",x"00001497",x"00001495",x"00001493",x"00001491",
		x"0000148f",x"0000148d",x"0000148b",x"00001489",x"00001487",x"00001485",x"00001483",x"00001481",
		x"0000147f",x"0000147d",x"0000147b",x"00001479",x"00001477",x"00001475",x"00001473",x"00001471",
		x"0000146f",x"0000146d",x"0000146b",x"00001469",x"00001467",x"00001465",x"00001463",x"00001461",
		x"0000145f",x"0000145d",x"0000145b",x"00001459",x"00001457",x"00001455",x"00001453",x"00001451",
		x"0000144f",x"0000144d",x"0000144b",x"00001449",x"00001447",x"00001445",x"00001443",x"00001441",
		x"0000143f",x"0000143d",x"0000143b",x"00001439",x"00001437",x"00001435",x"00001433",x"00001431",
		x"0000142f",x"0000142d",x"0000142b",x"00001429",x"00001427",x"00001425",x"00001423",x"00001421",
		x"0000141f",x"0000141d",x"0000141b",x"00001419",x"00001417",x"00001415",x"00001413",x"00001411",
		x"0000140f",x"0000140d",x"0000140b",x"00001409",x"00001407",x"00001405",x"00001403",x"00001401",
		x"000013ff",x"000013fd",x"000013fb",x"000013f9",x"000013f7",x"000013f5",x"000013f3",x"000013f1",
		x"000013ef",x"000013ed",x"000013eb",x"000013e9",x"000013e7",x"000013e5",x"000013e3",x"000013e1",
		x"000013df",x"000013dd",x"000013db",x"000013d9",x"000013d7",x"000013d5",x"000013d3",x"000013d1",
		x"000013cf",x"000013cd",x"000013cb",x"000013c9",x"000013c7",x"000013c5",x"000013c3",x"000013c1",
		x"000013bf",x"000013bd",x"000013bb",x"000013b9",x"000013b7",x"000013b5",x"000013b3",x"000013b1",
		x"000013af",x"000013ad",x"000013ab",x"000013a9",x"000013a7",x"000013a5",x"000013a3",x"000013a1",
		x"0000139f",x"0000139d",x"0000139b",x"00001399",x"00001397",x"00001395",x"00001393",x"00001391",
		x"0000138f",x"0000138d",x"0000138b",x"00001389",x"00001386",x"00001384",x"00001382",x"00001380",
		x"0000137e",x"0000137c",x"0000137a",x"00001378",x"00001376",x"00001374",x"00001372",x"00001370",
		x"0000136e",x"0000136c",x"0000136a",x"00001368",x"00001366",x"00001364",x"00001362",x"00001360",
		x"0000135e",x"0000135c",x"0000135a",x"00001358",x"00001356",x"00001354",x"00001352",x"00001350",
		x"0000134e",x"0000134c",x"0000134a",x"00001348",x"00001346",x"00001344",x"00001342",x"00001340",
		x"0000133e",x"0000133c",x"0000133a",x"00001338",x"00001336",x"00001334",x"00001332",x"00001330",
		x"0000132e",x"0000132c",x"0000132a",x"00001328",x"00001326",x"00001324",x"00001322",x"00001320",
		x"0000131e",x"0000131c",x"0000131a",x"00001318",x"00001316",x"00001314",x"00001312",x"00001310",
		x"0000130e",x"0000130c",x"0000130a",x"00001308",x"00001306",x"00001304",x"00001302",x"00001300",
		x"000012fe",x"000012fc",x"000012fa",x"000012f8",x"000012f6",x"000012f4",x"000012f2",x"000012f0",
		x"000012ee",x"000012ec",x"000012ea",x"000012e8",x"000012e6",x"000012e4",x"000012e2",x"000012e0",
		x"000012de",x"000012dc",x"000012da",x"000012d8",x"000012d6",x"000012d4",x"000012d2",x"000012d0",
		x"000012ce",x"000012cc",x"000012ca",x"000012c8",x"000012c6",x"000012c4",x"000012c2",x"000012c0",
		x"000012be",x"000012bc",x"000012ba",x"000012b8",x"000012b6",x"000012b4",x"000012b2",x"000012b0",
		x"000012ae",x"000012ac",x"000012aa",x"000012a8",x"000012a6",x"000012a4",x"000012a2",x"000012a0",
		x"0000129e",x"0000129c",x"0000129a",x"00001298",x"00001296",x"00001294",x"00001292",x"00001290",
		x"0000128e",x"0000128c",x"0000128a",x"00001288",x"00001286",x"00001284",x"00001282",x"00001280",
		x"0000127e",x"0000127c",x"0000127a",x"00001278",x"00001276",x"00001274",x"00001272",x"00001270",
		x"0000126e",x"0000126c",x"0000126a",x"00001268",x"00001266",x"00001264",x"00001262",x"00001260",
		x"0000125e",x"0000125c",x"0000125a",x"00001258",x"00001256",x"00001254",x"00001252",x"00001250",
		x"0000124e",x"0000124c",x"0000124a",x"00001248",x"00001246",x"00001244",x"00001242",x"00001240",
		x"0000123e",x"0000123c",x"0000123a",x"00001238",x"00001236",x"00001234",x"00001232",x"00001230",
		x"0000122e",x"0000122c",x"0000122a",x"00001228",x"00001226",x"00001224",x"00001222",x"00001220",
		x"0000121e",x"0000121c",x"0000121a",x"00001218",x"00001216",x"00001214",x"00001212",x"00001210",
		x"0000120e",x"0000120c",x"0000120a",x"00001208",x"00001206",x"00001204",x"00001202",x"00001200",
		x"000011fe",x"000011fc",x"000011fa",x"000011f8",x"000011f6",x"000011f4",x"000011f2",x"000011f0",
		x"000011ee",x"000011ec",x"000011ea",x"000011e8",x"000011e6",x"000011e4",x"000011e2",x"000011e0",
		x"000011de",x"000011dc",x"000011da",x"000011d8",x"000011d6",x"000011d4",x"000011d2",x"000011d0",
		x"000011ce",x"000011cc",x"000011ca",x"000011c8",x"000011c6",x"000011c4",x"000011c2",x"000011c0",
		x"000011be",x"000011bc",x"000011ba",x"000011b8",x"000011b6",x"000011b4",x"000011b2",x"000011b0",
		x"000011ae",x"000011ac",x"000011aa",x"000011a8",x"000011a6",x"000011a4",x"000011a2",x"000011a0",
		x"0000119e",x"0000119c",x"0000119a",x"00001198",x"00001196",x"00001194",x"00001192",x"00001190",
		x"0000118e",x"0000118c",x"0000118a",x"00001188",x"00001186",x"00001184",x"00001182",x"00001180",
		x"0000117e",x"0000117c",x"0000117a",x"00001178",x"00001176",x"00001174",x"00001172",x"00001170",
		x"0000116e",x"0000116c",x"0000116a",x"00001168",x"00001166",x"00001164",x"00001162",x"00001160",
		x"0000115e",x"0000115c",x"0000115a",x"00001158",x"00001156",x"00001154",x"00001152",x"00001150",
		x"0000114e",x"0000114c",x"0000114a",x"00001148",x"00001146",x"00001144",x"00001142",x"00001140",
		x"0000113e",x"0000113c",x"0000113a",x"00001138",x"00001136",x"00001134",x"00001132",x"00001130",
		x"0000112e",x"0000112c",x"0000112a",x"00001128",x"00001126",x"00001124",x"00001122",x"00001120",
		x"0000111e",x"0000111c",x"0000111a",x"00001118",x"00001116",x"00001114",x"00001112",x"00001110",
		x"0000110e",x"0000110c",x"0000110a",x"00001108",x"00001106",x"00001104",x"00001102",x"00001100",
		x"000010fe",x"000010fc",x"000010fa",x"000010f8",x"000010f6",x"000010f4",x"000010f2",x"000010f0",
		x"000010ee",x"000010ec",x"000010ea",x"000010e8",x"000010e6",x"000010e4",x"000010e2",x"000010e0",
		x"000010de",x"000010dc",x"000010da",x"000010d8",x"000010d6",x"000010d4",x"000010d2",x"000010d0",
		x"000010ce",x"000010cc",x"000010ca",x"000010c8",x"000010c6",x"000010c4",x"000010c2",x"000010c0",
		x"000010be",x"000010bc",x"000010ba",x"000010b8",x"000010b6",x"000010b4",x"000010b2",x"000010b0",
		x"000010ae",x"000010ac",x"000010aa",x"000010a8",x"000010a6",x"000010a4",x"000010a2",x"000010a0",
		x"0000109e",x"0000109c",x"0000109a",x"00001098",x"00001096",x"00001094",x"00001092",x"00001090",
		x"0000108e",x"0000108c",x"0000108a",x"00001088",x"00001086",x"00001084",x"00001082",x"00001080",
		x"0000107e",x"0000107c",x"0000107a",x"00001078",x"00001076",x"00001074",x"00001072",x"00001070",
		x"0000106e",x"0000106c",x"0000106a",x"00001068",x"00001066",x"00001064",x"00001062",x"00001060",
		x"0000105e",x"0000105c",x"0000105a",x"00001058",x"00001056",x"00001054",x"00001052",x"00001050",
		x"0000104e",x"0000104c",x"0000104a",x"00001048",x"00001046",x"00001044",x"00001042",x"00001040",
		x"0000103e",x"0000103c",x"0000103a",x"00001038",x"00001036",x"00001034",x"00001032",x"00001030",
		x"0000102e",x"0000102c",x"0000102a",x"00001028",x"00001026",x"00001024",x"00001022",x"00001020",
		x"0000101e",x"0000101c",x"0000101a",x"00001018",x"00001016",x"00001014",x"00001012",x"00001010",
		x"0000100e",x"0000100c",x"0000100a",x"00001008",x"00001006",x"00001004",x"00001002",x"00001000",
		x"00000ffe",x"00000ffc",x"00000ffa",x"00000ff8",x"00000ff6",x"00000ff4",x"00000ff2",x"00000ff0",
		x"00000fee",x"00000fec",x"00000fea",x"00000fe8",x"00000fe6",x"00000fe4",x"00000fe2",x"00000fe0",
		x"00000fde",x"00000fdc",x"00000fda",x"00000fd8",x"00000fd6",x"00000fd4",x"00000fd2",x"00000fd0",
		x"00000fce",x"00000fcc",x"00000fca",x"00000fc8",x"00000fc6",x"00000fc4",x"00000fc2",x"00000fc0",
		x"00000fbe",x"00000fbc",x"00000fba",x"00000fb8",x"00000fb6",x"00000fb4",x"00000fb2",x"00000fb0",
		x"00000fae",x"00000fac",x"00000faa",x"00000fa8",x"00000fa6",x"00000fa4",x"00000fa2",x"00000fa0",
		x"00000f9e",x"00000f9c",x"00000f9a",x"00000f98",x"00000f96",x"00000f94",x"00000f92",x"00000f90",
		x"00000f8e",x"00000f8c",x"00000f8a",x"00000f88",x"00000f86",x"00000f84",x"00000f82",x"00000f80",
		x"00000f7e",x"00000f7c",x"00000f7a",x"00000f78",x"00000f76",x"00000f74",x"00000f72",x"00000f70",
		x"00000f6e",x"00000f6c",x"00000f6a",x"00000f68",x"00000f66",x"00000f64",x"00000f62",x"00000f60",
		x"00000f5e",x"00000f5c",x"00000f5a",x"00000f58",x"00000f56",x"00000f54",x"00000f52",x"00000f50",
		x"00000f4e",x"00000f4c",x"00000f4a",x"00000f48",x"00000f46",x"00000f44",x"00000f42",x"00000f40",
		x"00000f3e",x"00000f3c",x"00000f3a",x"00000f38",x"00000f36",x"00000f34",x"00000f32",x"00000f30",
		x"00000f2e",x"00000f2c",x"00000f2a",x"00000f28",x"00000f26",x"00000f24",x"00000f22",x"00000f20",
		x"00000f1e",x"00000f1c",x"00000f1a",x"00000f18",x"00000f16",x"00000f14",x"00000f12",x"00000f10",
		x"00000f0e",x"00000f0c",x"00000f0a",x"00000f08",x"00000f06",x"00000f04",x"00000f02",x"00000f00",
		x"00000efe",x"00000efc",x"00000efa",x"00000ef8",x"00000ef6",x"00000ef4",x"00000ef2",x"00000ef0",
		x"00000eee",x"00000eec",x"00000eea",x"00000ee8",x"00000ee6",x"00000ee4",x"00000ee2",x"00000ee0",
		x"00000ede",x"00000edc",x"00000eda",x"00000ed8",x"00000ed6",x"00000ed4",x"00000ed2",x"00000ed0",
		x"00000ece",x"00000ecc",x"00000eca",x"00000ec8",x"00000ec6",x"00000ec4",x"00000ec2",x"00000ec0",
		x"00000ebe",x"00000ebc",x"00000eba",x"00000eb8",x"00000eb6",x"00000eb4",x"00000eb2",x"00000eb0",
		x"00000eae",x"00000eac",x"00000eaa",x"00000ea8",x"00000ea6",x"00000ea4",x"00000ea2",x"00000ea0",
		x"00000e9e",x"00000e9c",x"00000e9a",x"00000e98",x"00000e96",x"00000e94",x"00000e92",x"00000e90",
		x"00000e8e",x"00000e8c",x"00000e8a",x"00000e88",x"00000e86",x"00000e84",x"00000e82",x"00000e80",
		x"00000e7e",x"00000e7c",x"00000e7a",x"00000e78",x"00000e76",x"00000e74",x"00000e72",x"00000e70",
		x"00000e6e",x"00000e6c",x"00000e6a",x"00000e68",x"00000e66",x"00000e64",x"00000e62",x"00000e60",
		x"00000e5e",x"00000e5c",x"00000e5a",x"00000e58",x"00000e56",x"00000e54",x"00000e52",x"00000e50",
		x"00000e4e",x"00000e4c",x"00000e4a",x"00000e48",x"00000e46",x"00000e44",x"00000e42",x"00000e40",
		x"00000e3e",x"00000e3c",x"00000e3a",x"00000e38",x"00000e36",x"00000e34",x"00000e32",x"00000e30",
		x"00000e2e",x"00000e2c",x"00000e2a",x"00000e28",x"00000e26",x"00000e24",x"00000e22",x"00000e20",
		x"00000e1e",x"00000e1c",x"00000e1a",x"00000e18",x"00000e16",x"00000e14",x"00000e12",x"00000e10",
		x"00000e0e",x"00000e0c",x"00000e0a",x"00000e08",x"00000e06",x"00000e04",x"00000e02",x"00000e00",
		x"00000dfe",x"00000dfc",x"00000dfa",x"00000df8",x"00000df6",x"00000df4",x"00000df2",x"00000df0",
		x"00000dee",x"00000dec",x"00000dea",x"00000de8",x"00000de6",x"00000de4",x"00000de2",x"00000de0",
		x"00000dde",x"00000ddc",x"00000dda",x"00000dd8",x"00000dd6",x"00000dd4",x"00000dd2",x"00000dd0",
		x"00000dce",x"00000dcc",x"00000dca",x"00000dc8",x"00000dc6",x"00000dc4",x"00000dc2",x"00000dc0",
		x"00000dbe",x"00000dbc",x"00000dba",x"00000db8",x"00000db6",x"00000db4",x"00000db2",x"00000db0",
		x"00000dae",x"00000dac",x"00000daa",x"00000da8",x"00000da6",x"00000da4",x"00000da2",x"00000da0",
		x"00000d9e",x"00000d9c",x"00000d9a",x"00000d98",x"00000d96",x"00000d94",x"00000d92",x"00000d90",
		x"00000d8e",x"00000d8c",x"00000d8a",x"00000d88",x"00000d86",x"00000d84",x"00000d82",x"00000d80",
		x"00000d7e",x"00000d7c",x"00000d7a",x"00000d78",x"00000d76",x"00000d74",x"00000d72",x"00000d70",
		x"00000d6e",x"00000d6c",x"00000d6a",x"00000d68",x"00000d66",x"00000d64",x"00000d62",x"00000d60",
		x"00000d5e",x"00000d5c",x"00000d5a",x"00000d58",x"00000d56",x"00000d54",x"00000d52",x"00000d50",
		x"00000d4e",x"00000d4c",x"00000d4a",x"00000d48",x"00000d46",x"00000d44",x"00000d42",x"00000d40",
		x"00000d3e",x"00000d3c",x"00000d3a",x"00000d38",x"00000d36",x"00000d34",x"00000d32",x"00000d30",
		x"00000d2e",x"00000d2c",x"00000d2a",x"00000d28",x"00000d26",x"00000d24",x"00000d22",x"00000d20",
		x"00000d1e",x"00000d1c",x"00000d1a",x"00000d18",x"00000d16",x"00000d14",x"00000d12",x"00000d10",
		x"00000d0e",x"00000d0c",x"00000d0a",x"00000d08",x"00000d06",x"00000d04",x"00000d02",x"00000d00",
		x"00000cfe",x"00000cfc",x"00000cfa",x"00000cf8",x"00000cf6",x"00000cf4",x"00000cf2",x"00000cf0",
		x"00000cee",x"00000cec",x"00000cea",x"00000ce8",x"00000ce6",x"00000ce4",x"00000ce2",x"00000ce0",
		x"00000cde",x"00000cdc",x"00000cda",x"00000cd8",x"00000cd6",x"00000cd4",x"00000cd2",x"00000cd0",
		x"00000cce",x"00000ccc",x"00000cca",x"00000cc8",x"00000cc6",x"00000cc4",x"00000cc2",x"00000cc0",
		x"00000cbe",x"00000cbc",x"00000cba",x"00000cb8",x"00000cb6",x"00000cb4",x"00000cb2",x"00000cb0",
		x"00000cae",x"00000cac",x"00000caa",x"00000ca8",x"00000ca6",x"00000ca4",x"00000ca2",x"00000ca0",
		x"00000c9e",x"00000c9c",x"00000c9a",x"00000c98",x"00000c96",x"00000c94",x"00000c92",x"00000c90",
		x"00000c8e",x"00000c8c",x"00000c8a",x"00000c88",x"00000c86",x"00000c84",x"00000c82",x"00000c80",
		x"00000c7e",x"00000c7c",x"00000c7a",x"00000c78",x"00000c76",x"00000c74",x"00000c72",x"00000c70",
		x"00000c6e",x"00000c6c",x"00000c6a",x"00000c68",x"00000c66",x"00000c64",x"00000c62",x"00000c60",
		x"00000c5e",x"00000c5c",x"00000c5a",x"00000c58",x"00000c56",x"00000c54",x"00000c52",x"00000c50",
		x"00000c4e",x"00000c4c",x"00000c4a",x"00000c48",x"00000c46",x"00000c44",x"00000c42",x"00000c40",
		x"00000c3e",x"00000c3c",x"00000c3a",x"00000c38",x"00000c36",x"00000c34",x"00000c32",x"00000c30",
		x"00000c2e",x"00000c2c",x"00000c2a",x"00000c28",x"00000c26",x"00000c24",x"00000c22",x"00000c20",
		x"00000c1e",x"00000c1c",x"00000c1a",x"00000c18",x"00000c16",x"00000c14",x"00000c12",x"00000c10",
		x"00000c0e",x"00000c0c",x"00000c0a",x"00000c08",x"00000c06",x"00000c04",x"00000c02",x"00000c00",
		x"00000bfe",x"00000bfc",x"00000bfa",x"00000bf8",x"00000bf6",x"00000bf4",x"00000bf2",x"00000bf0",
		x"00000bee",x"00000bec",x"00000bea",x"00000be8",x"00000be6",x"00000be4",x"00000be2",x"00000be0",
		x"00000bde",x"00000bdc",x"00000bda",x"00000bd8",x"00000bd6",x"00000bd4",x"00000bd2",x"00000bd0",
		x"00000bce",x"00000bcc",x"00000bca",x"00000bc8",x"00000bc6",x"00000bc4",x"00000bc2",x"00000bc0",
		x"00000bbe",x"00000bbc",x"00000bba",x"00000bb8",x"00000bb6",x"00000bb4",x"00000bb2",x"00000bb0",
		x"00000bae",x"00000bac",x"00000baa",x"00000ba8",x"00000ba6",x"00000ba4",x"00000ba2",x"00000ba0",
		x"00000b9e",x"00000b9c",x"00000b9a",x"00000b98",x"00000b96",x"00000b94",x"00000b92",x"00000b90",
		x"00000b8e",x"00000b8c",x"00000b8a",x"00000b88",x"00000b86",x"00000b84",x"00000b82",x"00000b80",
		x"00000b7e",x"00000b7c",x"00000b7a",x"00000b78",x"00000b76",x"00000b74",x"00000b72",x"00000b70",
		x"00000b6e",x"00000b6c",x"00000b6a",x"00000b68",x"00000b66",x"00000b64",x"00000b62",x"00000b60",
		x"00000b5e",x"00000b5c",x"00000b5a",x"00000b58",x"00000b56",x"00000b54",x"00000b52",x"00000b50",
		x"00000b4e",x"00000b4c",x"00000b4a",x"00000b48",x"00000b46",x"00000b44",x"00000b42",x"00000b40",
		x"00000b3e",x"00000b3c",x"00000b3a",x"00000b38",x"00000b36",x"00000b34",x"00000b32",x"00000b30",
		x"00000b2e",x"00000b2c",x"00000b2a",x"00000b28",x"00000b26",x"00000b24",x"00000b22",x"00000b20",
		x"00000b1e",x"00000b1c",x"00000b1a",x"00000b18",x"00000b16",x"00000b14",x"00000b12",x"00000b10",
		x"00000b0e",x"00000b0c",x"00000b0a",x"00000b08",x"00000b06",x"00000b04",x"00000b02",x"00000b00",
		x"00000afe",x"00000afc",x"00000afa",x"00000af8",x"00000af6",x"00000af4",x"00000af2",x"00000af0",
		x"00000aee",x"00000aec",x"00000aea",x"00000ae8",x"00000ae6",x"00000ae4",x"00000ae2",x"00000ae0",
		x"00000ade",x"00000adc",x"00000ada",x"00000ad8",x"00000ad6",x"00000ad4",x"00000ad2",x"00000ad0",
		x"00000ace",x"00000acc",x"00000aca",x"00000ac8",x"00000ac6",x"00000ac4",x"00000ac2",x"00000ac0",
		x"00000abe",x"00000abc",x"00000aba",x"00000ab8",x"00000ab6",x"00000ab4",x"00000ab2",x"00000ab0",
		x"00000aae",x"00000aac",x"00000aaa",x"00000aa8",x"00000aa6",x"00000aa4",x"00000aa2",x"00000aa0",
		x"00000a9e",x"00000a9c",x"00000a9a",x"00000a98",x"00000a96",x"00000a94",x"00000a92",x"00000a90",
		x"00000a8e",x"00000a8c",x"00000a8a",x"00000a88",x"00000a86",x"00000a84",x"00000a82",x"00000a80",
		x"00000a7e",x"00000a7c",x"00000a7a",x"00000a78",x"00000a76",x"00000a74",x"00000a72",x"00000a70",
		x"00000a6e",x"00000a6c",x"00000a6a",x"00000a68",x"00000a66",x"00000a64",x"00000a62",x"00000a60",
		x"00000a5e",x"00000a5c",x"00000a5a",x"00000a58",x"00000a56",x"00000a54",x"00000a52",x"00000a50",
		x"00000a4e",x"00000a4c",x"00000a4a",x"00000a48",x"00000a46",x"00000a44",x"00000a42",x"00000a40",
		x"00000a3e",x"00000a3c",x"00000a3a",x"00000a38",x"00000a36",x"00000a34",x"00000a32",x"00000a30",
		x"00000a2e",x"00000a2c",x"00000a2a",x"00000a28",x"00000a26",x"00000a24",x"00000a22",x"00000a20",
		x"00000a1e",x"00000a1c",x"00000a1a",x"00000a18",x"00000a16",x"00000a14",x"00000a12",x"00000a10",
		x"00000a0e",x"00000a0c",x"00000a0a",x"00000a08",x"00000a06",x"00000a04",x"00000a02",x"00000a00",
		x"000009fe",x"000009fc",x"000009fa",x"000009f8",x"000009f6",x"000009f4",x"000009f2",x"000009f0",
		x"000009ee",x"000009ec",x"000009ea",x"000009e8",x"000009e6",x"000009e4",x"000009e2",x"000009e0",
		x"000009de",x"000009dc",x"000009da",x"000009d8",x"000009d6",x"000009d4",x"000009d2",x"000009d0",
		x"000009ce",x"000009cc",x"000009ca",x"000009c8",x"000009c6",x"000009c4",x"000009c2",x"000009c0",
		x"000009be",x"000009bc",x"000009ba",x"000009b8",x"000009b6",x"000009b4",x"000009b2",x"000009b0",
		x"000009ae",x"000009ac",x"000009aa",x"000009a8",x"000009a6",x"000009a4",x"000009a2",x"000009a0",
		x"0000099e",x"0000099c",x"0000099a",x"00000998",x"00000996",x"00000994",x"00000992",x"00000990",
		x"0000098e",x"0000098c",x"0000098a",x"00000988",x"00000986",x"00000984",x"00000982",x"00000980",
		x"0000097e",x"0000097c",x"0000097a",x"00000978",x"00000976",x"00000974",x"00000972",x"00000970",
		x"0000096e",x"0000096c",x"0000096a",x"00000968",x"00000966",x"00000964",x"00000962",x"00000960",
		x"0000095e",x"0000095c",x"0000095a",x"00000958",x"00000956",x"00000954",x"00000952",x"00000950",
		x"0000094e",x"0000094c",x"0000094a",x"00000948",x"00000946",x"00000944",x"00000942",x"00000940",
		x"0000093e",x"0000093c",x"0000093a",x"00000938",x"00000936",x"00000934",x"00000932",x"00000930",
		x"0000092e",x"0000092c",x"0000092a",x"00000928",x"00000926",x"00000924",x"00000922",x"00000920",
		x"0000091e",x"0000091c",x"0000091a",x"00000918",x"00000916",x"00000914",x"00000912",x"00000910",
		x"0000090e",x"0000090c",x"0000090a",x"00000908",x"00000906",x"00000904",x"00000902",x"00000900",
		x"000008fe",x"000008fc",x"000008fa",x"000008f8",x"000008f6",x"000008f4",x"000008f2",x"000008f0",
		x"000008ee",x"000008ec",x"000008ea",x"000008e8",x"000008e6",x"000008e4",x"000008e2",x"000008e0",
		x"000008de",x"000008dc",x"000008da",x"000008d8",x"000008d6",x"000008d4",x"000008d2",x"000008d0",
		x"000008ce",x"000008cc",x"000008ca",x"000008c8",x"000008c6",x"000008c4",x"000008c2",x"000008c0",
		x"000008be",x"000008bc",x"000008ba",x"000008b8",x"000008b6",x"000008b4",x"000008b2",x"000008b0",
		x"000008ae",x"000008ac",x"000008aa",x"000008a8",x"000008a6",x"000008a4",x"000008a2",x"000008a0",
		x"0000089e",x"0000089c",x"0000089a",x"00000898",x"00000896",x"00000894",x"00000892",x"00000890",
		x"0000088e",x"0000088c",x"0000088a",x"00000888",x"00000886",x"00000884",x"00000882",x"00000880",
		x"0000087e",x"0000087c",x"0000087a",x"00000878",x"00000876",x"00000874",x"00000872",x"00000870",
		x"0000086e",x"0000086c",x"0000086a",x"00000868",x"00000866",x"00000864",x"00000862",x"00000860",
		x"0000085e",x"0000085c",x"0000085a",x"00000858",x"00000856",x"00000854",x"00000852",x"00000850",
		x"0000084e",x"0000084c",x"0000084a",x"00000848",x"00000846",x"00000844",x"00000842",x"00000840",
		x"0000083e",x"0000083c",x"0000083a",x"00000838",x"00000836",x"00000834",x"00000832",x"00000830",
		x"0000082e",x"0000082c",x"0000082a",x"00000828",x"00000826",x"00000824",x"00000822",x"00000820",
		x"0000081e",x"0000081c",x"0000081a",x"00000818",x"00000816",x"00000814",x"00000812",x"00000810",
		x"0000080e",x"0000080c",x"0000080a",x"00000808",x"00000806",x"00000804",x"00000802",x"00000800",
		x"000007fe",x"000007fc",x"000007fa",x"000007f8",x"000007f6",x"000007f4",x"000007f2",x"000007f0",
		x"000007ee",x"000007ec",x"000007ea",x"000007e8",x"000007e6",x"000007e4",x"000007e2",x"000007e0",
		x"000007de",x"000007dc",x"000007da",x"000007d8",x"000007d6",x"000007d4",x"000007d2",x"000007d0",
		x"000007ce",x"000007cc",x"000007ca",x"000007c8",x"000007c6",x"000007c4",x"000007c2",x"000007c0",
		x"000007be",x"000007bc",x"000007ba",x"000007b8",x"000007b6",x"000007b4",x"000007b2",x"000007b0",
		x"000007ae",x"000007ac",x"000007aa",x"000007a8",x"000007a6",x"000007a4",x"000007a2",x"000007a0",
		x"0000079e",x"0000079c",x"0000079a",x"00000798",x"00000796",x"00000794",x"00000792",x"00000790",
		x"0000078e",x"0000078c",x"0000078a",x"00000788",x"00000786",x"00000784",x"00000782",x"00000780",
		x"0000077e",x"0000077c",x"0000077a",x"00000778",x"00000776",x"00000774",x"00000772",x"00000770",
		x"0000076e",x"0000076c",x"0000076a",x"00000768",x"00000766",x"00000764",x"00000762",x"00000760",
		x"0000075e",x"0000075c",x"0000075a",x"00000758",x"00000756",x"00000754",x"00000752",x"00000750",
		x"0000074e",x"0000074c",x"0000074a",x"00000748",x"00000746",x"00000744",x"00000742",x"00000740",
		x"0000073e",x"0000073c",x"0000073a",x"00000738",x"00000736",x"00000734",x"00000732",x"00000730",
		x"0000072e",x"0000072c",x"0000072a",x"00000728",x"00000726",x"00000724",x"00000722",x"00000720",
		x"0000071e",x"0000071c",x"0000071a",x"00000718",x"00000716",x"00000714",x"00000712",x"00000710",
		x"0000070e",x"0000070c",x"0000070a",x"00000708",x"00000706",x"00000704",x"00000702",x"00000700",
		x"000006fe",x"000006fc",x"000006fa",x"000006f8",x"000006f6",x"000006f4",x"000006f2",x"000006f0",
		x"000006ee",x"000006ec",x"000006ea",x"000006e8",x"000006e6",x"000006e4",x"000006e2",x"000006e0",
		x"000006de",x"000006dc",x"000006da",x"000006d8",x"000006d6",x"000006d4",x"000006d2",x"000006d0",
		x"000006ce",x"000006cc",x"000006ca",x"000006c8",x"000006c6",x"000006c4",x"000006c2",x"000006c0",
		x"000006be",x"000006bc",x"000006ba",x"000006b8",x"000006b6",x"000006b4",x"000006b2",x"000006b0",
		x"000006ae",x"000006ac",x"000006aa",x"000006a8",x"000006a6",x"000006a4",x"000006a2",x"000006a0",
		x"0000069e",x"0000069c",x"0000069a",x"00000698",x"00000696",x"00000694",x"00000692",x"00000690",
		x"0000068e",x"0000068c",x"0000068a",x"00000688",x"00000686",x"00000684",x"00000682",x"00000680",
		x"0000067e",x"0000067c",x"0000067a",x"00000678",x"00000676",x"00000674",x"00000672",x"00000670",
		x"0000066e",x"0000066c",x"0000066a",x"00000668",x"00000666",x"00000664",x"00000662",x"00000660",
		x"0000065e",x"0000065c",x"0000065a",x"00000658",x"00000656",x"00000654",x"00000652",x"00000650",
		x"0000064e",x"0000064c",x"0000064a",x"00000648",x"00000646",x"00000644",x"00000642",x"00000640",
		x"0000063e",x"0000063c",x"0000063a",x"00000638",x"00000636",x"00000634",x"00000632",x"00000630",
		x"0000062e",x"0000062c",x"0000062a",x"00000628",x"00000626",x"00000624",x"00000622",x"00000620",
		x"0000061e",x"0000061c",x"0000061a",x"00000618",x"00000616",x"00000614",x"00000612",x"00000610",
		x"0000060e",x"0000060c",x"0000060a",x"00000608",x"00000606",x"00000604",x"00000602",x"00000600",
		x"000005fe",x"000005fc",x"000005fa",x"000005f8",x"000005f6",x"000005f4",x"000005f2",x"000005f0",
		x"000005ee",x"000005ec",x"000005ea",x"000005e8",x"000005e6",x"000005e4",x"000005e2",x"000005e0",
		x"000005de",x"000005dc",x"000005da",x"000005d8",x"000005d6",x"000005d4",x"000005d2",x"000005d0",
		x"000005ce",x"000005cc",x"000005ca",x"000005c8",x"000005c6",x"000005c4",x"000005c2",x"000005c0",
		x"000005be",x"000005bc",x"000005ba",x"000005b8",x"000005b6",x"000005b4",x"000005b2",x"000005b0",
		x"000005ae",x"000005ac",x"000005aa",x"000005a8",x"000005a6",x"000005a4",x"000005a2",x"000005a0",
		x"0000059e",x"0000059c",x"0000059a",x"00000598",x"00000596",x"00000594",x"00000592",x"00000590",
		x"0000058e",x"0000058c",x"0000058a",x"00000588",x"00000586",x"00000584",x"00000582",x"00000580",
		x"0000057e",x"0000057c",x"0000057a",x"00000578",x"00000576",x"00000574",x"00000572",x"00000570",
		x"0000056e",x"0000056c",x"0000056a",x"00000568",x"00000566",x"00000564",x"00000562",x"00000560",
		x"0000055e",x"0000055c",x"0000055a",x"00000558",x"00000556",x"00000554",x"00000552",x"00000550",
		x"0000054e",x"0000054c",x"0000054a",x"00000548",x"00000546",x"00000544",x"00000542",x"00000540",
		x"0000053e",x"0000053c",x"0000053a",x"00000538",x"00000536",x"00000534",x"00000532",x"00000530",
		x"0000052e",x"0000052c",x"0000052a",x"00000528",x"00000526",x"00000524",x"00000522",x"00000520",
		x"0000051e",x"0000051c",x"0000051a",x"00000518",x"00000516",x"00000514",x"00000512",x"00000510",
		x"0000050e",x"0000050c",x"0000050a",x"00000508",x"00000506",x"00000504",x"00000502",x"00000500",
		x"000004fe",x"000004fc",x"000004fa",x"000004f8",x"000004f6",x"000004f4",x"000004f2",x"000004f0",
		x"000004ee",x"000004ec",x"000004ea",x"000004e8",x"000004e6",x"000004e4",x"000004e2",x"000004e0",
		x"000004de",x"000004dc",x"000004da",x"000004d8",x"000004d6",x"000004d4",x"000004d2",x"000004d0",
		x"000004ce",x"000004cc",x"000004ca",x"000004c8",x"000004c6",x"000004c4",x"000004c2",x"000004c0",
		x"000004be",x"000004bc",x"000004ba",x"000004b8",x"000004b6",x"000004b4",x"000004b2",x"000004b0",
		x"000004ae",x"000004ac",x"000004aa",x"000004a8",x"000004a6",x"000004a4",x"000004a2",x"000004a0",
		x"0000049e",x"0000049c",x"0000049a",x"00000498",x"00000496",x"00000494",x"00000492",x"00000490",
		x"0000048e",x"0000048c",x"0000048a",x"00000488",x"00000486",x"00000484",x"00000482",x"00000480",
		x"0000047e",x"0000047c",x"0000047a",x"00000478",x"00000476",x"00000474",x"00000472",x"00000470",
		x"0000046e",x"0000046c",x"0000046a",x"00000468",x"00000466",x"00000464",x"00000462",x"00000460",
		x"0000045e",x"0000045c",x"0000045a",x"00000458",x"00000456",x"00000454",x"00000452",x"00000450",
		x"0000044e",x"0000044c",x"0000044a",x"00000448",x"00000446",x"00000444",x"00000442",x"00000440",
		x"0000043e",x"0000043c",x"0000043a",x"00000438",x"00000436",x"00000434",x"00000432",x"00000430",
		x"0000042e",x"0000042c",x"0000042a",x"00000428",x"00000426",x"00000424",x"00000422",x"00000420",
		x"0000041e",x"0000041c",x"0000041a",x"00000418",x"00000416",x"00000414",x"00000412",x"00000410",
		x"0000040e",x"0000040c",x"0000040a",x"00000408",x"00000406",x"00000404",x"00000402",x"00000400",
		x"000003fe",x"000003fc",x"000003fa",x"000003f8",x"000003f6",x"000003f4",x"000003f2",x"000003f0",
		x"000003ee",x"000003ec",x"000003ea",x"000003e8",x"000003e6",x"000003e4",x"000003e2",x"000003e0",
		x"000003de",x"000003dc",x"000003da",x"000003d8",x"000003d6",x"000003d4",x"000003d2",x"000003d0",
		x"000003ce",x"000003cc",x"000003ca",x"000003c8",x"000003c6",x"000003c4",x"000003c2",x"000003c0",
		x"000003be",x"000003bc",x"000003ba",x"000003b8",x"000003b6",x"000003b4",x"000003b2",x"000003b0",
		x"000003ae",x"000003ac",x"000003aa",x"000003a8",x"000003a6",x"000003a4",x"000003a2",x"000003a0",
		x"0000039e",x"0000039c",x"0000039a",x"00000398",x"00000396",x"00000394",x"00000392",x"00000390",
		x"0000038e",x"0000038c",x"0000038a",x"00000388",x"00000386",x"00000384",x"00000382",x"00000380",
		x"0000037e",x"0000037c",x"0000037a",x"00000378",x"00000376",x"00000374",x"00000372",x"00000370",
		x"0000036e",x"0000036c",x"0000036a",x"00000368",x"00000366",x"00000364",x"00000362",x"00000360",
		x"0000035e",x"0000035c",x"0000035a",x"00000358",x"00000356",x"00000354",x"00000352",x"00000350",
		x"0000034e",x"0000034c",x"0000034a",x"00000348",x"00000346",x"00000344",x"00000342",x"00000340",
		x"0000033e",x"0000033c",x"0000033a",x"00000338",x"00000336",x"00000334",x"00000332",x"00000330",
		x"0000032e",x"0000032c",x"0000032a",x"00000328",x"00000326",x"00000324",x"00000322",x"00000320",
		x"0000031e",x"0000031c",x"0000031a",x"00000318",x"00000316",x"00000314",x"00000312",x"00000310",
		x"0000030e",x"0000030c",x"0000030a",x"00000308",x"00000306",x"00000304",x"00000302",x"00000300",
		x"000002fe",x"000002fc",x"000002fa",x"000002f8",x"000002f6",x"000002f4",x"000002f2",x"000002f0",
		x"000002ee",x"000002ec",x"000002ea",x"000002e8",x"000002e6",x"000002e4",x"000002e2",x"000002e0",
		x"000002de",x"000002dc",x"000002da",x"000002d8",x"000002d6",x"000002d4",x"000002d2",x"000002d0",
		x"000002ce",x"000002cc",x"000002ca",x"000002c8",x"000002c6",x"000002c4",x"000002c2",x"000002c0",
		x"000002be",x"000002bc",x"000002ba",x"000002b8",x"000002b6",x"000002b4",x"000002b2",x"000002b0",
		x"000002ae",x"000002ac",x"000002aa",x"000002a8",x"000002a6",x"000002a4",x"000002a2",x"000002a0",
		x"0000029e",x"0000029c",x"0000029a",x"00000298",x"00000296",x"00000294",x"00000292",x"00000290",
		x"0000028e",x"0000028c",x"0000028a",x"00000288",x"00000286",x"00000284",x"00000282",x"00000280",
		x"0000027e",x"0000027c",x"0000027a",x"00000278",x"00000276",x"00000274",x"00000272",x"00000270",
		x"0000026e",x"0000026c",x"0000026a",x"00000268",x"00000266",x"00000264",x"00000262",x"00000260",
		x"0000025e",x"0000025c",x"0000025a",x"00000258",x"00000256",x"00000254",x"00000252",x"00000250",
		x"0000024e",x"0000024c",x"0000024a",x"00000248",x"00000246",x"00000244",x"00000242",x"00000240",
		x"0000023e",x"0000023c",x"0000023a",x"00000238",x"00000236",x"00000234",x"00000232",x"00000230",
		x"0000022e",x"0000022c",x"0000022a",x"00000228",x"00000226",x"00000224",x"00000222",x"00000220",
		x"0000021e",x"0000021c",x"0000021a",x"00000218",x"00000216",x"00000214",x"00000212",x"00000210",
		x"0000020e",x"0000020c",x"0000020a",x"00000208",x"00000206",x"00000204",x"00000202",x"00000200",
		x"000001fe",x"000001fc",x"000001fa",x"000001f8",x"000001f6",x"000001f4",x"000001f2",x"000001f0",
		x"000001ee",x"000001ec",x"000001ea",x"000001e8",x"000001e6",x"000001e4",x"000001e2",x"000001e0",
		x"000001de",x"000001dc",x"000001da",x"000001d8",x"000001d6",x"000001d4",x"000001d2",x"000001d0",
		x"000001ce",x"000001cc",x"000001ca",x"000001c8",x"000001c6",x"000001c4",x"000001c2",x"000001c0",
		x"000001be",x"000001bc",x"000001ba",x"000001b8",x"000001b6",x"000001b4",x"000001b2",x"000001b0",
		x"000001ae",x"000001ac",x"000001aa",x"000001a8",x"000001a6",x"000001a4",x"000001a2",x"000001a0",
		x"0000019e",x"0000019c",x"0000019a",x"00000198",x"00000196",x"00000194",x"00000192",x"00000190",
		x"0000018e",x"0000018c",x"0000018a",x"00000188",x"00000186",x"00000184",x"00000182",x"00000180",
		x"0000017e",x"0000017c",x"0000017a",x"00000178",x"00000176",x"00000174",x"00000172",x"00000170",
		x"0000016e",x"0000016c",x"0000016a",x"00000168",x"00000166",x"00000164",x"00000162",x"00000160",
		x"0000015e",x"0000015c",x"0000015a",x"00000158",x"00000156",x"00000154",x"00000152",x"00000150",
		x"0000014e",x"0000014c",x"0000014a",x"00000148",x"00000146",x"00000144",x"00000142",x"00000140",
		x"0000013e",x"0000013c",x"0000013a",x"00000138",x"00000136",x"00000134",x"00000132",x"00000130",
		x"0000012e",x"0000012c",x"0000012a",x"00000128",x"00000126",x"00000124",x"00000122",x"00000120",
		x"0000011e",x"0000011c",x"0000011a",x"00000118",x"00000116",x"00000114",x"00000112",x"00000110",
		x"0000010e",x"0000010c",x"0000010a",x"00000108",x"00000106",x"00000104",x"00000102",x"00000100",
		x"000000fe",x"000000fc",x"000000fa",x"000000f8",x"000000f6",x"000000f4",x"000000f2",x"000000f0",
		x"000000ee",x"000000ec",x"000000ea",x"000000e8",x"000000e6",x"000000e4",x"000000e2",x"000000e0",
		x"000000de",x"000000dc",x"000000da",x"000000d8",x"000000d6",x"000000d4",x"000000d2",x"000000d0",
		x"000000ce",x"000000cc",x"000000ca",x"000000c8",x"000000c6",x"000000c4",x"000000c2",x"000000c0",
		x"000000be",x"000000bc",x"000000ba",x"000000b8",x"000000b6",x"000000b4",x"000000b2",x"000000b0",
		x"000000ae",x"000000ac",x"000000aa",x"000000a8",x"000000a6",x"000000a4",x"000000a2",x"000000a0",
		x"0000009e",x"0000009c",x"0000009a",x"00000098",x"00000096",x"00000094",x"00000092",x"00000090",
		x"0000008e",x"0000008c",x"0000008a",x"00000088",x"00000086",x"00000084",x"00000082",x"00000080",
		x"0000007e",x"0000007c",x"0000007a",x"00000078",x"00000076",x"00000074",x"00000072",x"00000070",
		x"0000006e",x"0000006c",x"0000006a",x"00000068",x"00000066",x"00000064",x"00000062",x"00000060",
		x"0000005e",x"0000005c",x"0000005a",x"00000058",x"00000056",x"00000054",x"00000052",x"00000050",
		x"0000004e",x"0000004c",x"0000004a",x"00000048",x"00000046",x"00000044",x"00000042",x"00000040",
		x"0000003e",x"0000003c",x"0000003a",x"00000038",x"00000036",x"00000034",x"00000032",x"00000030",
		x"0000002e",x"0000002c",x"0000002a",x"00000028",x"00000026",x"00000024",x"00000022",x"00000020",
		x"0000001e",x"0000001c",x"0000001a",x"00000018",x"00000016",x"00000014",x"00000012",x"00000010",
		x"0000000e",x"0000000c",x"0000000a",x"00000008",x"00000006",x"00000004",x"00000002",x"00000000"
	);
begin
    
	process (clk)
		variable counter:	std_logic_vector(32-1 downto 0) := (others => '0');
		variable index: integer range 1 to 10001 := 1;
		--variable cociente : std_logic_vector(32-1 downto 0) := (others => '0');
		variable cociente : integer range 1 to 60000 :=1;
		variable resto : integer range 0 to 60000 :=0;
	begin
		if (rising_edge(clk)) then
			counter := counter + 10000;--antes era 100.
			-- if counter >= 1000  =  10ns * 1000 = 10 000ns
			--    increment index and reset counter
--			if (counter >= frq) then
--				index := index + 1;
--				counter:=counter-frq;
--				while(counter>frq)loop
--					index := index + 1;
--					counter:=counter-frq;
--				end loop;
--				--counter := (others => '0');
--			end if;

			if (counter >= frq) then
				cociente:=((to_integer(unsigned(std_logic_vector(counter))))/(to_integer(unsigned(std_logic_vector(frq)))));
				index:=index + cociente;
				resto:=((to_integer(unsigned(std_logic_vector(counter))))rem(to_integer(unsigned(std_logic_vector(frq)))));
				counter:= std_logic_vector(to_unsigned(resto, 32));
				--counter := (others => '0');
			end if;

			-- if index > 100 reset it to 1
			if (index > 10000) then
				index := 1;
			end if;
		end if;
		pwm_ctrl <= data(index);
	end process;

end Behavioral;
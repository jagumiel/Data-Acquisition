library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use ieee.numeric_std.all;
--use ieee.numeric_std;


entity sin is
	port (
		clk:		in	std_logic;
		amp:		in	std_logic_vector(32-1 downto 0);--La puedes quitar.
		frq:		in	std_logic_vector(32-1 downto 0);
		pwm_ctrl:	out	std_logic_vector(32-1 downto 0)
	);
end sin;

architecture Behavioral of sin is

	type  SAMPLE_main is array (1 to 10000) of std_logic_vector(31 downto 0);
	constant data : SAMPLE_main := (
		x"00001388",x"0000138b",x"0000138e",x"00001391",x"00001395",x"00001398",x"0000139b",x"0000139e",
		x"000013a1",x"000013a4",x"000013a7",x"000013ab",x"000013ae",x"000013b1",x"000013b4",x"000013b7",
		x"000013ba",x"000013bd",x"000013c1",x"000013c4",x"000013c7",x"000013ca",x"000013cd",x"000013d0",
		x"000013d3",x"000013d7",x"000013da",x"000013dd",x"000013e0",x"000013e3",x"000013e6",x"000013e9",
		x"000013ed",x"000013f0",x"000013f3",x"000013f6",x"000013f9",x"000013fc",x"000013ff",x"00001403",
		x"00001406",x"00001409",x"0000140c",x"0000140f",x"00001412",x"00001415",x"00001419",x"0000141c",
		x"0000141f",x"00001422",x"00001425",x"00001428",x"0000142b",x"0000142e",x"00001432",x"00001435",
		x"00001438",x"0000143b",x"0000143e",x"00001441",x"00001444",x"00001448",x"0000144b",x"0000144e",
		x"00001451",x"00001454",x"00001457",x"0000145a",x"0000145e",x"00001461",x"00001464",x"00001467",
		x"0000146a",x"0000146d",x"00001470",x"00001474",x"00001477",x"0000147a",x"0000147d",x"00001480",
		x"00001483",x"00001486",x"0000148a",x"0000148d",x"00001490",x"00001493",x"00001496",x"00001499",
		x"0000149c",x"0000149f",x"000014a3",x"000014a6",x"000014a9",x"000014ac",x"000014af",x"000014b2",
		x"000014b5",x"000014b9",x"000014bc",x"000014bf",x"000014c2",x"000014c5",x"000014c8",x"000014cb",
		x"000014cf",x"000014d2",x"000014d5",x"000014d8",x"000014db",x"000014de",x"000014e1",x"000014e4",
		x"000014e8",x"000014eb",x"000014ee",x"000014f1",x"000014f4",x"000014f7",x"000014fa",x"000014fe",
		x"00001501",x"00001504",x"00001507",x"0000150a",x"0000150d",x"00001510",x"00001513",x"00001517",
		x"0000151a",x"0000151d",x"00001520",x"00001523",x"00001526",x"00001529",x"0000152d",x"00001530",
		x"00001533",x"00001536",x"00001539",x"0000153c",x"0000153f",x"00001542",x"00001546",x"00001549",
		x"0000154c",x"0000154f",x"00001552",x"00001555",x"00001558",x"0000155b",x"0000155f",x"00001562",
		x"00001565",x"00001568",x"0000156b",x"0000156e",x"00001571",x"00001574",x"00001578",x"0000157b",
		x"0000157e",x"00001581",x"00001584",x"00001587",x"0000158a",x"0000158d",x"00001591",x"00001594",
		x"00001597",x"0000159a",x"0000159d",x"000015a0",x"000015a3",x"000015a6",x"000015aa",x"000015ad",
		x"000015b0",x"000015b3",x"000015b6",x"000015b9",x"000015bc",x"000015bf",x"000015c3",x"000015c6",
		x"000015c9",x"000015cc",x"000015cf",x"000015d2",x"000015d5",x"000015d8",x"000015dc",x"000015df",
		x"000015e2",x"000015e5",x"000015e8",x"000015eb",x"000015ee",x"000015f1",x"000015f4",x"000015f8",
		x"000015fb",x"000015fe",x"00001601",x"00001604",x"00001607",x"0000160a",x"0000160d",x"00001611",
		x"00001614",x"00001617",x"0000161a",x"0000161d",x"00001620",x"00001623",x"00001626",x"00001629",
		x"0000162d",x"00001630",x"00001633",x"00001636",x"00001639",x"0000163c",x"0000163f",x"00001642",
		x"00001645",x"00001649",x"0000164c",x"0000164f",x"00001652",x"00001655",x"00001658",x"0000165b",
		x"0000165e",x"00001661",x"00001665",x"00001668",x"0000166b",x"0000166e",x"00001671",x"00001674",
		x"00001677",x"0000167a",x"0000167d",x"00001681",x"00001684",x"00001687",x"0000168a",x"0000168d",
		x"00001690",x"00001693",x"00001696",x"00001699",x"0000169c",x"000016a0",x"000016a3",x"000016a6",
		x"000016a9",x"000016ac",x"000016af",x"000016b2",x"000016b5",x"000016b8",x"000016bb",x"000016bf",
		x"000016c2",x"000016c5",x"000016c8",x"000016cb",x"000016ce",x"000016d1",x"000016d4",x"000016d7",
		x"000016da",x"000016de",x"000016e1",x"000016e4",x"000016e7",x"000016ea",x"000016ed",x"000016f0",
		x"000016f3",x"000016f6",x"000016f9",x"000016fc",x"00001700",x"00001703",x"00001706",x"00001709",
		x"0000170c",x"0000170f",x"00001712",x"00001715",x"00001718",x"0000171b",x"0000171e",x"00001722",
		x"00001725",x"00001728",x"0000172b",x"0000172e",x"00001731",x"00001734",x"00001737",x"0000173a",
		x"0000173d",x"00001740",x"00001744",x"00001747",x"0000174a",x"0000174d",x"00001750",x"00001753",
		x"00001756",x"00001759",x"0000175c",x"0000175f",x"00001762",x"00001765",x"00001768",x"0000176c",
		x"0000176f",x"00001772",x"00001775",x"00001778",x"0000177b",x"0000177e",x"00001781",x"00001784",
		x"00001787",x"0000178a",x"0000178d",x"00001790",x"00001794",x"00001797",x"0000179a",x"0000179d",
		x"000017a0",x"000017a3",x"000017a6",x"000017a9",x"000017ac",x"000017af",x"000017b2",x"000017b5",
		x"000017b8",x"000017bb",x"000017bf",x"000017c2",x"000017c5",x"000017c8",x"000017cb",x"000017ce",
		x"000017d1",x"000017d4",x"000017d7",x"000017da",x"000017dd",x"000017e0",x"000017e3",x"000017e6",
		x"000017e9",x"000017ed",x"000017f0",x"000017f3",x"000017f6",x"000017f9",x"000017fc",x"000017ff",
		x"00001802",x"00001805",x"00001808",x"0000180b",x"0000180e",x"00001811",x"00001814",x"00001817",
		x"0000181a",x"0000181d",x"00001821",x"00001824",x"00001827",x"0000182a",x"0000182d",x"00001830",
		x"00001833",x"00001836",x"00001839",x"0000183c",x"0000183f",x"00001842",x"00001845",x"00001848",
		x"0000184b",x"0000184e",x"00001851",x"00001854",x"00001857",x"0000185a",x"0000185d",x"00001861",
		x"00001864",x"00001867",x"0000186a",x"0000186d",x"00001870",x"00001873",x"00001876",x"00001879",
		x"0000187c",x"0000187f",x"00001882",x"00001885",x"00001888",x"0000188b",x"0000188e",x"00001891",
		x"00001894",x"00001897",x"0000189a",x"0000189d",x"000018a0",x"000018a3",x"000018a6",x"000018a9",
		x"000018ac",x"000018af",x"000018b3",x"000018b6",x"000018b9",x"000018bc",x"000018bf",x"000018c2",
		x"000018c5",x"000018c8",x"000018cb",x"000018ce",x"000018d1",x"000018d4",x"000018d7",x"000018da",
		x"000018dd",x"000018e0",x"000018e3",x"000018e6",x"000018e9",x"000018ec",x"000018ef",x"000018f2",
		x"000018f5",x"000018f8",x"000018fb",x"000018fe",x"00001901",x"00001904",x"00001907",x"0000190a",
		x"0000190d",x"00001910",x"00001913",x"00001916",x"00001919",x"0000191c",x"0000191f",x"00001922",
		x"00001925",x"00001928",x"0000192b",x"0000192e",x"00001931",x"00001934",x"00001937",x"0000193a",
		x"0000193d",x"00001940",x"00001943",x"00001946",x"00001949",x"0000194c",x"0000194f",x"00001952",
		x"00001955",x"00001958",x"0000195b",x"0000195e",x"00001961",x"00001964",x"00001967",x"0000196a",
		x"0000196d",x"00001970",x"00001973",x"00001976",x"00001979",x"0000197c",x"0000197f",x"00001982",
		x"00001985",x"00001988",x"0000198b",x"0000198e",x"00001991",x"00001994",x"00001997",x"0000199a",
		x"0000199d",x"000019a0",x"000019a3",x"000019a6",x"000019a9",x"000019ac",x"000019af",x"000019b2",
		x"000019b5",x"000019b8",x"000019bb",x"000019be",x"000019c1",x"000019c4",x"000019c7",x"000019ca",
		x"000019cd",x"000019d0",x"000019d3",x"000019d6",x"000019d9",x"000019dc",x"000019df",x"000019e2",
		x"000019e5",x"000019e8",x"000019eb",x"000019ee",x"000019f1",x"000019f4",x"000019f6",x"000019f9",
		x"000019fc",x"000019ff",x"00001a02",x"00001a05",x"00001a08",x"00001a0b",x"00001a0e",x"00001a11",
		x"00001a14",x"00001a17",x"00001a1a",x"00001a1d",x"00001a20",x"00001a23",x"00001a26",x"00001a29",
		x"00001a2c",x"00001a2f",x"00001a32",x"00001a35",x"00001a38",x"00001a3b",x"00001a3d",x"00001a40",
		x"00001a43",x"00001a46",x"00001a49",x"00001a4c",x"00001a4f",x"00001a52",x"00001a55",x"00001a58",
		x"00001a5b",x"00001a5e",x"00001a61",x"00001a64",x"00001a67",x"00001a6a",x"00001a6d",x"00001a70",
		x"00001a72",x"00001a75",x"00001a78",x"00001a7b",x"00001a7e",x"00001a81",x"00001a84",x"00001a87",
		x"00001a8a",x"00001a8d",x"00001a90",x"00001a93",x"00001a96",x"00001a99",x"00001a9c",x"00001a9e",
		x"00001aa1",x"00001aa4",x"00001aa7",x"00001aaa",x"00001aad",x"00001ab0",x"00001ab3",x"00001ab6",
		x"00001ab9",x"00001abc",x"00001abf",x"00001ac2",x"00001ac4",x"00001ac7",x"00001aca",x"00001acd",
		x"00001ad0",x"00001ad3",x"00001ad6",x"00001ad9",x"00001adc",x"00001adf",x"00001ae2",x"00001ae5",
		x"00001ae7",x"00001aea",x"00001aed",x"00001af0",x"00001af3",x"00001af6",x"00001af9",x"00001afc",
		x"00001aff",x"00001b02",x"00001b05",x"00001b07",x"00001b0a",x"00001b0d",x"00001b10",x"00001b13",
		x"00001b16",x"00001b19",x"00001b1c",x"00001b1f",x"00001b21",x"00001b24",x"00001b27",x"00001b2a",
		x"00001b2d",x"00001b30",x"00001b33",x"00001b36",x"00001b39",x"00001b3b",x"00001b3e",x"00001b41",
		x"00001b44",x"00001b47",x"00001b4a",x"00001b4d",x"00001b50",x"00001b53",x"00001b55",x"00001b58",
		x"00001b5b",x"00001b5e",x"00001b61",x"00001b64",x"00001b67",x"00001b6a",x"00001b6c",x"00001b6f",
		x"00001b72",x"00001b75",x"00001b78",x"00001b7b",x"00001b7e",x"00001b81",x"00001b83",x"00001b86",
		x"00001b89",x"00001b8c",x"00001b8f",x"00001b92",x"00001b95",x"00001b97",x"00001b9a",x"00001b9d",
		x"00001ba0",x"00001ba3",x"00001ba6",x"00001ba9",x"00001bac",x"00001bae",x"00001bb1",x"00001bb4",
		x"00001bb7",x"00001bba",x"00001bbd",x"00001bbf",x"00001bc2",x"00001bc5",x"00001bc8",x"00001bcb",
		x"00001bce",x"00001bd1",x"00001bd3",x"00001bd6",x"00001bd9",x"00001bdc",x"00001bdf",x"00001be2",
		x"00001be4",x"00001be7",x"00001bea",x"00001bed",x"00001bf0",x"00001bf3",x"00001bf5",x"00001bf8",
		x"00001bfb",x"00001bfe",x"00001c01",x"00001c04",x"00001c06",x"00001c09",x"00001c0c",x"00001c0f",
		x"00001c12",x"00001c15",x"00001c17",x"00001c1a",x"00001c1d",x"00001c20",x"00001c23",x"00001c26",
		x"00001c28",x"00001c2b",x"00001c2e",x"00001c31",x"00001c34",x"00001c36",x"00001c39",x"00001c3c",
		x"00001c3f",x"00001c42",x"00001c45",x"00001c47",x"00001c4a",x"00001c4d",x"00001c50",x"00001c53",
		x"00001c55",x"00001c58",x"00001c5b",x"00001c5e",x"00001c61",x"00001c63",x"00001c66",x"00001c69",
		x"00001c6c",x"00001c6f",x"00001c71",x"00001c74",x"00001c77",x"00001c7a",x"00001c7d",x"00001c7f",
		x"00001c82",x"00001c85",x"00001c88",x"00001c8a",x"00001c8d",x"00001c90",x"00001c93",x"00001c96",
		x"00001c98",x"00001c9b",x"00001c9e",x"00001ca1",x"00001ca4",x"00001ca6",x"00001ca9",x"00001cac",
		x"00001caf",x"00001cb1",x"00001cb4",x"00001cb7",x"00001cba",x"00001cbd",x"00001cbf",x"00001cc2",
		x"00001cc5",x"00001cc8",x"00001cca",x"00001ccd",x"00001cd0",x"00001cd3",x"00001cd5",x"00001cd8",
		x"00001cdb",x"00001cde",x"00001ce0",x"00001ce3",x"00001ce6",x"00001ce9",x"00001ceb",x"00001cee",
		x"00001cf1",x"00001cf4",x"00001cf6",x"00001cf9",x"00001cfc",x"00001cff",x"00001d01",x"00001d04",
		x"00001d07",x"00001d0a",x"00001d0c",x"00001d0f",x"00001d12",x"00001d15",x"00001d17",x"00001d1a",
		x"00001d1d",x"00001d20",x"00001d22",x"00001d25",x"00001d28",x"00001d2b",x"00001d2d",x"00001d30",
		x"00001d33",x"00001d36",x"00001d38",x"00001d3b",x"00001d3e",x"00001d40",x"00001d43",x"00001d46",
		x"00001d49",x"00001d4b",x"00001d4e",x"00001d51",x"00001d53",x"00001d56",x"00001d59",x"00001d5c",
		x"00001d5e",x"00001d61",x"00001d64",x"00001d66",x"00001d69",x"00001d6c",x"00001d6f",x"00001d71",
		x"00001d74",x"00001d77",x"00001d79",x"00001d7c",x"00001d7f",x"00001d82",x"00001d84",x"00001d87",
		x"00001d8a",x"00001d8c",x"00001d8f",x"00001d92",x"00001d94",x"00001d97",x"00001d9a",x"00001d9d",
		x"00001d9f",x"00001da2",x"00001da5",x"00001da7",x"00001daa",x"00001dad",x"00001daf",x"00001db2",
		x"00001db5",x"00001db7",x"00001dba",x"00001dbd",x"00001dbf",x"00001dc2",x"00001dc5",x"00001dc7",
		x"00001dca",x"00001dcd",x"00001dcf",x"00001dd2",x"00001dd5",x"00001dd7",x"00001dda",x"00001ddd",
		x"00001ddf",x"00001de2",x"00001de5",x"00001de7",x"00001dea",x"00001ded",x"00001def",x"00001df2",
		x"00001df5",x"00001df7",x"00001dfa",x"00001dfd",x"00001dff",x"00001e02",x"00001e05",x"00001e07",
		x"00001e0a",x"00001e0d",x"00001e0f",x"00001e12",x"00001e15",x"00001e17",x"00001e1a",x"00001e1c",
		x"00001e1f",x"00001e22",x"00001e24",x"00001e27",x"00001e2a",x"00001e2c",x"00001e2f",x"00001e32",
		x"00001e34",x"00001e37",x"00001e39",x"00001e3c",x"00001e3f",x"00001e41",x"00001e44",x"00001e47",
		x"00001e49",x"00001e4c",x"00001e4e",x"00001e51",x"00001e54",x"00001e56",x"00001e59",x"00001e5c",
		x"00001e5e",x"00001e61",x"00001e63",x"00001e66",x"00001e69",x"00001e6b",x"00001e6e",x"00001e70",
		x"00001e73",x"00001e76",x"00001e78",x"00001e7b",x"00001e7d",x"00001e80",x"00001e83",x"00001e85",
		x"00001e88",x"00001e8a",x"00001e8d",x"00001e90",x"00001e92",x"00001e95",x"00001e97",x"00001e9a",
		x"00001e9d",x"00001e9f",x"00001ea2",x"00001ea4",x"00001ea7",x"00001eaa",x"00001eac",x"00001eaf",
		x"00001eb1",x"00001eb4",x"00001eb6",x"00001eb9",x"00001ebc",x"00001ebe",x"00001ec1",x"00001ec3",
		x"00001ec6",x"00001ec8",x"00001ecb",x"00001ece",x"00001ed0",x"00001ed3",x"00001ed5",x"00001ed8",
		x"00001eda",x"00001edd",x"00001edf",x"00001ee2",x"00001ee5",x"00001ee7",x"00001eea",x"00001eec",
		x"00001eef",x"00001ef1",x"00001ef4",x"00001ef6",x"00001ef9",x"00001efc",x"00001efe",x"00001f01",
		x"00001f03",x"00001f06",x"00001f08",x"00001f0b",x"00001f0d",x"00001f10",x"00001f12",x"00001f15",
		x"00001f17",x"00001f1a",x"00001f1d",x"00001f1f",x"00001f22",x"00001f24",x"00001f27",x"00001f29",
		x"00001f2c",x"00001f2e",x"00001f31",x"00001f33",x"00001f36",x"00001f38",x"00001f3b",x"00001f3d",
		x"00001f40",x"00001f42",x"00001f45",x"00001f47",x"00001f4a",x"00001f4c",x"00001f4f",x"00001f51",
		x"00001f54",x"00001f56",x"00001f59",x"00001f5b",x"00001f5e",x"00001f60",x"00001f63",x"00001f65",
		x"00001f68",x"00001f6a",x"00001f6d",x"00001f6f",x"00001f72",x"00001f74",x"00001f77",x"00001f79",
		x"00001f7c",x"00001f7e",x"00001f81",x"00001f83",x"00001f86",x"00001f88",x"00001f8b",x"00001f8d",
		x"00001f90",x"00001f92",x"00001f95",x"00001f97",x"00001f9a",x"00001f9c",x"00001f9e",x"00001fa1",
		x"00001fa3",x"00001fa6",x"00001fa8",x"00001fab",x"00001fad",x"00001fb0",x"00001fb2",x"00001fb5",
		x"00001fb7",x"00001fba",x"00001fbc",x"00001fbe",x"00001fc1",x"00001fc3",x"00001fc6",x"00001fc8",
		x"00001fcb",x"00001fcd",x"00001fd0",x"00001fd2",x"00001fd4",x"00001fd7",x"00001fd9",x"00001fdc",
		x"00001fde",x"00001fe1",x"00001fe3",x"00001fe6",x"00001fe8",x"00001fea",x"00001fed",x"00001fef",
		x"00001ff2",x"00001ff4",x"00001ff7",x"00001ff9",x"00001ffb",x"00001ffe",x"00002000",x"00002003",
		x"00002005",x"00002007",x"0000200a",x"0000200c",x"0000200f",x"00002011",x"00002014",x"00002016",
		x"00002018",x"0000201b",x"0000201d",x"00002020",x"00002022",x"00002024",x"00002027",x"00002029",
		x"0000202c",x"0000202e",x"00002030",x"00002033",x"00002035",x"00002038",x"0000203a",x"0000203c",
		x"0000203f",x"00002041",x"00002043",x"00002046",x"00002048",x"0000204b",x"0000204d",x"0000204f",
		x"00002052",x"00002054",x"00002056",x"00002059",x"0000205b",x"0000205e",x"00002060",x"00002062",
		x"00002065",x"00002067",x"00002069",x"0000206c",x"0000206e",x"00002070",x"00002073",x"00002075",
		x"00002078",x"0000207a",x"0000207c",x"0000207f",x"00002081",x"00002083",x"00002086",x"00002088",
		x"0000208a",x"0000208d",x"0000208f",x"00002091",x"00002094",x"00002096",x"00002098",x"0000209b",
		x"0000209d",x"0000209f",x"000020a2",x"000020a4",x"000020a6",x"000020a9",x"000020ab",x"000020ad",
		x"000020b0",x"000020b2",x"000020b4",x"000020b7",x"000020b9",x"000020bb",x"000020be",x"000020c0",
		x"000020c2",x"000020c5",x"000020c7",x"000020c9",x"000020cb",x"000020ce",x"000020d0",x"000020d2",
		x"000020d5",x"000020d7",x"000020d9",x"000020dc",x"000020de",x"000020e0",x"000020e2",x"000020e5",
		x"000020e7",x"000020e9",x"000020ec",x"000020ee",x"000020f0",x"000020f2",x"000020f5",x"000020f7",
		x"000020f9",x"000020fc",x"000020fe",x"00002100",x"00002102",x"00002105",x"00002107",x"00002109",
		x"0000210b",x"0000210e",x"00002110",x"00002112",x"00002115",x"00002117",x"00002119",x"0000211b",
		x"0000211e",x"00002120",x"00002122",x"00002124",x"00002127",x"00002129",x"0000212b",x"0000212d",
		x"00002130",x"00002132",x"00002134",x"00002136",x"00002139",x"0000213b",x"0000213d",x"0000213f",
		x"00002142",x"00002144",x"00002146",x"00002148",x"0000214a",x"0000214d",x"0000214f",x"00002151",
		x"00002153",x"00002156",x"00002158",x"0000215a",x"0000215c",x"0000215e",x"00002161",x"00002163",
		x"00002165",x"00002167",x"0000216a",x"0000216c",x"0000216e",x"00002170",x"00002172",x"00002175",
		x"00002177",x"00002179",x"0000217b",x"0000217d",x"00002180",x"00002182",x"00002184",x"00002186",
		x"00002188",x"0000218b",x"0000218d",x"0000218f",x"00002191",x"00002193",x"00002195",x"00002198",
		x"0000219a",x"0000219c",x"0000219e",x"000021a0",x"000021a3",x"000021a5",x"000021a7",x"000021a9",
		x"000021ab",x"000021ad",x"000021b0",x"000021b2",x"000021b4",x"000021b6",x"000021b8",x"000021ba",
		x"000021bd",x"000021bf",x"000021c1",x"000021c3",x"000021c5",x"000021c7",x"000021c9",x"000021cc",
		x"000021ce",x"000021d0",x"000021d2",x"000021d4",x"000021d6",x"000021d8",x"000021db",x"000021dd",
		x"000021df",x"000021e1",x"000021e3",x"000021e5",x"000021e7",x"000021e9",x"000021ec",x"000021ee",
		x"000021f0",x"000021f2",x"000021f4",x"000021f6",x"000021f8",x"000021fa",x"000021fd",x"000021ff",
		x"00002201",x"00002203",x"00002205",x"00002207",x"00002209",x"0000220b",x"0000220d",x"00002210",
		x"00002212",x"00002214",x"00002216",x"00002218",x"0000221a",x"0000221c",x"0000221e",x"00002220",
		x"00002222",x"00002224",x"00002227",x"00002229",x"0000222b",x"0000222d",x"0000222f",x"00002231",
		x"00002233",x"00002235",x"00002237",x"00002239",x"0000223b",x"0000223d",x"0000223f",x"00002241",
		x"00002244",x"00002246",x"00002248",x"0000224a",x"0000224c",x"0000224e",x"00002250",x"00002252",
		x"00002254",x"00002256",x"00002258",x"0000225a",x"0000225c",x"0000225e",x"00002260",x"00002262",
		x"00002264",x"00002266",x"00002268",x"0000226a",x"0000226c",x"0000226f",x"00002271",x"00002273",
		x"00002275",x"00002277",x"00002279",x"0000227b",x"0000227d",x"0000227f",x"00002281",x"00002283",
		x"00002285",x"00002287",x"00002289",x"0000228b",x"0000228d",x"0000228f",x"00002291",x"00002293",
		x"00002295",x"00002297",x"00002299",x"0000229b",x"0000229d",x"0000229f",x"000022a1",x"000022a3",
		x"000022a5",x"000022a7",x"000022a9",x"000022ab",x"000022ad",x"000022af",x"000022b1",x"000022b3",
		x"000022b5",x"000022b7",x"000022b9",x"000022bb",x"000022bd",x"000022bf",x"000022c1",x"000022c3",
		x"000022c4",x"000022c6",x"000022c8",x"000022ca",x"000022cc",x"000022ce",x"000022d0",x"000022d2",
		x"000022d4",x"000022d6",x"000022d8",x"000022da",x"000022dc",x"000022de",x"000022e0",x"000022e2",
		x"000022e4",x"000022e6",x"000022e8",x"000022ea",x"000022eb",x"000022ed",x"000022ef",x"000022f1",
		x"000022f3",x"000022f5",x"000022f7",x"000022f9",x"000022fb",x"000022fd",x"000022ff",x"00002301",
		x"00002303",x"00002304",x"00002306",x"00002308",x"0000230a",x"0000230c",x"0000230e",x"00002310",
		x"00002312",x"00002314",x"00002316",x"00002318",x"00002319",x"0000231b",x"0000231d",x"0000231f",
		x"00002321",x"00002323",x"00002325",x"00002327",x"00002329",x"0000232a",x"0000232c",x"0000232e",
		x"00002330",x"00002332",x"00002334",x"00002336",x"00002338",x"00002339",x"0000233b",x"0000233d",
		x"0000233f",x"00002341",x"00002343",x"00002345",x"00002347",x"00002348",x"0000234a",x"0000234c",
		x"0000234e",x"00002350",x"00002352",x"00002354",x"00002355",x"00002357",x"00002359",x"0000235b",
		x"0000235d",x"0000235f",x"00002360",x"00002362",x"00002364",x"00002366",x"00002368",x"0000236a",
		x"0000236b",x"0000236d",x"0000236f",x"00002371",x"00002373",x"00002375",x"00002376",x"00002378",
		x"0000237a",x"0000237c",x"0000237e",x"0000237f",x"00002381",x"00002383",x"00002385",x"00002387",
		x"00002388",x"0000238a",x"0000238c",x"0000238e",x"00002390",x"00002391",x"00002393",x"00002395",
		x"00002397",x"00002399",x"0000239a",x"0000239c",x"0000239e",x"000023a0",x"000023a1",x"000023a3",
		x"000023a5",x"000023a7",x"000023a9",x"000023aa",x"000023ac",x"000023ae",x"000023b0",x"000023b1",
		x"000023b3",x"000023b5",x"000023b7",x"000023b8",x"000023ba",x"000023bc",x"000023be",x"000023c0",
		x"000023c1",x"000023c3",x"000023c5",x"000023c6",x"000023c8",x"000023ca",x"000023cc",x"000023cd",
		x"000023cf",x"000023d1",x"000023d3",x"000023d4",x"000023d6",x"000023d8",x"000023da",x"000023db",
		x"000023dd",x"000023df",x"000023e0",x"000023e2",x"000023e4",x"000023e6",x"000023e7",x"000023e9",
		x"000023eb",x"000023ec",x"000023ee",x"000023f0",x"000023f2",x"000023f3",x"000023f5",x"000023f7",
		x"000023f8",x"000023fa",x"000023fc",x"000023fd",x"000023ff",x"00002401",x"00002403",x"00002404",
		x"00002406",x"00002408",x"00002409",x"0000240b",x"0000240d",x"0000240e",x"00002410",x"00002412",
		x"00002413",x"00002415",x"00002417",x"00002418",x"0000241a",x"0000241c",x"0000241d",x"0000241f",
		x"00002421",x"00002422",x"00002424",x"00002426",x"00002427",x"00002429",x"0000242b",x"0000242c",
		x"0000242e",x"0000242f",x"00002431",x"00002433",x"00002434",x"00002436",x"00002438",x"00002439",
		x"0000243b",x"0000243d",x"0000243e",x"00002440",x"00002441",x"00002443",x"00002445",x"00002446",
		x"00002448",x"0000244a",x"0000244b",x"0000244d",x"0000244e",x"00002450",x"00002452",x"00002453",
		x"00002455",x"00002456",x"00002458",x"0000245a",x"0000245b",x"0000245d",x"0000245e",x"00002460",
		x"00002462",x"00002463",x"00002465",x"00002466",x"00002468",x"00002469",x"0000246b",x"0000246d",
		x"0000246e",x"00002470",x"00002471",x"00002473",x"00002474",x"00002476",x"00002478",x"00002479",
		x"0000247b",x"0000247c",x"0000247e",x"0000247f",x"00002481",x"00002483",x"00002484",x"00002486",
		x"00002487",x"00002489",x"0000248a",x"0000248c",x"0000248d",x"0000248f",x"00002490",x"00002492",
		x"00002494",x"00002495",x"00002497",x"00002498",x"0000249a",x"0000249b",x"0000249d",x"0000249e",
		x"000024a0",x"000024a1",x"000024a3",x"000024a4",x"000024a6",x"000024a7",x"000024a9",x"000024aa",
		x"000024ac",x"000024ad",x"000024af",x"000024b0",x"000024b2",x"000024b3",x"000024b5",x"000024b6",
		x"000024b8",x"000024b9",x"000024bb",x"000024bc",x"000024be",x"000024bf",x"000024c1",x"000024c2",
		x"000024c4",x"000024c5",x"000024c7",x"000024c8",x"000024ca",x"000024cb",x"000024cd",x"000024ce",
		x"000024cf",x"000024d1",x"000024d2",x"000024d4",x"000024d5",x"000024d7",x"000024d8",x"000024da",
		x"000024db",x"000024dd",x"000024de",x"000024df",x"000024e1",x"000024e2",x"000024e4",x"000024e5",
		x"000024e7",x"000024e8",x"000024ea",x"000024eb",x"000024ec",x"000024ee",x"000024ef",x"000024f1",
		x"000024f2",x"000024f4",x"000024f5",x"000024f6",x"000024f8",x"000024f9",x"000024fb",x"000024fc",
		x"000024fd",x"000024ff",x"00002500",x"00002502",x"00002503",x"00002504",x"00002506",x"00002507",
		x"00002509",x"0000250a",x"0000250b",x"0000250d",x"0000250e",x"00002510",x"00002511",x"00002512",
		x"00002514",x"00002515",x"00002517",x"00002518",x"00002519",x"0000251b",x"0000251c",x"0000251d",
		x"0000251f",x"00002520",x"00002521",x"00002523",x"00002524",x"00002526",x"00002527",x"00002528",
		x"0000252a",x"0000252b",x"0000252c",x"0000252e",x"0000252f",x"00002530",x"00002532",x"00002533",
		x"00002534",x"00002536",x"00002537",x"00002538",x"0000253a",x"0000253b",x"0000253c",x"0000253e",
		x"0000253f",x"00002540",x"00002542",x"00002543",x"00002544",x"00002546",x"00002547",x"00002548",
		x"0000254a",x"0000254b",x"0000254c",x"0000254d",x"0000254f",x"00002550",x"00002551",x"00002553",
		x"00002554",x"00002555",x"00002557",x"00002558",x"00002559",x"0000255a",x"0000255c",x"0000255d",
		x"0000255e",x"00002560",x"00002561",x"00002562",x"00002563",x"00002565",x"00002566",x"00002567",
		x"00002568",x"0000256a",x"0000256b",x"0000256c",x"0000256d",x"0000256f",x"00002570",x"00002571",
		x"00002573",x"00002574",x"00002575",x"00002576",x"00002577",x"00002579",x"0000257a",x"0000257b",
		x"0000257c",x"0000257e",x"0000257f",x"00002580",x"00002581",x"00002583",x"00002584",x"00002585",
		x"00002586",x"00002588",x"00002589",x"0000258a",x"0000258b",x"0000258c",x"0000258e",x"0000258f",
		x"00002590",x"00002591",x"00002592",x"00002594",x"00002595",x"00002596",x"00002597",x"00002598",
		x"0000259a",x"0000259b",x"0000259c",x"0000259d",x"0000259e",x"000025a0",x"000025a1",x"000025a2",
		x"000025a3",x"000025a4",x"000025a5",x"000025a7",x"000025a8",x"000025a9",x"000025aa",x"000025ab",
		x"000025ac",x"000025ae",x"000025af",x"000025b0",x"000025b1",x"000025b2",x"000025b3",x"000025b5",
		x"000025b6",x"000025b7",x"000025b8",x"000025b9",x"000025ba",x"000025bb",x"000025bd",x"000025be",
		x"000025bf",x"000025c0",x"000025c1",x"000025c2",x"000025c3",x"000025c4",x"000025c6",x"000025c7",
		x"000025c8",x"000025c9",x"000025ca",x"000025cb",x"000025cc",x"000025cd",x"000025cf",x"000025d0",
		x"000025d1",x"000025d2",x"000025d3",x"000025d4",x"000025d5",x"000025d6",x"000025d7",x"000025d8",
		x"000025da",x"000025db",x"000025dc",x"000025dd",x"000025de",x"000025df",x"000025e0",x"000025e1",
		x"000025e2",x"000025e3",x"000025e4",x"000025e5",x"000025e6",x"000025e8",x"000025e9",x"000025ea",
		x"000025eb",x"000025ec",x"000025ed",x"000025ee",x"000025ef",x"000025f0",x"000025f1",x"000025f2",
		x"000025f3",x"000025f4",x"000025f5",x"000025f6",x"000025f7",x"000025f8",x"000025f9",x"000025fa",
		x"000025fb",x"000025fc",x"000025fe",x"000025ff",x"00002600",x"00002601",x"00002602",x"00002603",
		x"00002604",x"00002605",x"00002606",x"00002607",x"00002608",x"00002609",x"0000260a",x"0000260b",
		x"0000260c",x"0000260d",x"0000260e",x"0000260f",x"00002610",x"00002611",x"00002612",x"00002613",
		x"00002614",x"00002615",x"00002616",x"00002617",x"00002618",x"00002619",x"0000261a",x"0000261b",
		x"0000261b",x"0000261c",x"0000261d",x"0000261e",x"0000261f",x"00002620",x"00002621",x"00002622",
		x"00002623",x"00002624",x"00002625",x"00002626",x"00002627",x"00002628",x"00002629",x"0000262a",
		x"0000262b",x"0000262c",x"0000262d",x"0000262e",x"0000262f",x"0000262f",x"00002630",x"00002631",
		x"00002632",x"00002633",x"00002634",x"00002635",x"00002636",x"00002637",x"00002638",x"00002639",
		x"0000263a",x"0000263a",x"0000263b",x"0000263c",x"0000263d",x"0000263e",x"0000263f",x"00002640",
		x"00002641",x"00002642",x"00002643",x"00002643",x"00002644",x"00002645",x"00002646",x"00002647",
		x"00002648",x"00002649",x"0000264a",x"0000264b",x"0000264b",x"0000264c",x"0000264d",x"0000264e",
		x"0000264f",x"00002650",x"00002651",x"00002651",x"00002652",x"00002653",x"00002654",x"00002655",
		x"00002656",x"00002657",x"00002657",x"00002658",x"00002659",x"0000265a",x"0000265b",x"0000265c",
		x"0000265c",x"0000265d",x"0000265e",x"0000265f",x"00002660",x"00002661",x"00002661",x"00002662",
		x"00002663",x"00002664",x"00002665",x"00002666",x"00002666",x"00002667",x"00002668",x"00002669",
		x"0000266a",x"0000266a",x"0000266b",x"0000266c",x"0000266d",x"0000266e",x"0000266e",x"0000266f",
		x"00002670",x"00002671",x"00002672",x"00002672",x"00002673",x"00002674",x"00002675",x"00002675",
		x"00002676",x"00002677",x"00002678",x"00002678",x"00002679",x"0000267a",x"0000267b",x"0000267c",
		x"0000267c",x"0000267d",x"0000267e",x"0000267f",x"0000267f",x"00002680",x"00002681",x"00002682",
		x"00002682",x"00002683",x"00002684",x"00002685",x"00002685",x"00002686",x"00002687",x"00002687",
		x"00002688",x"00002689",x"0000268a",x"0000268a",x"0000268b",x"0000268c",x"0000268d",x"0000268d",
		x"0000268e",x"0000268f",x"0000268f",x"00002690",x"00002691",x"00002691",x"00002692",x"00002693",
		x"00002694",x"00002694",x"00002695",x"00002696",x"00002696",x"00002697",x"00002698",x"00002698",
		x"00002699",x"0000269a",x"0000269a",x"0000269b",x"0000269c",x"0000269c",x"0000269d",x"0000269e",
		x"0000269e",x"0000269f",x"000026a0",x"000026a0",x"000026a1",x"000026a2",x"000026a2",x"000026a3",
		x"000026a4",x"000026a4",x"000026a5",x"000026a6",x"000026a6",x"000026a7",x"000026a8",x"000026a8",
		x"000026a9",x"000026aa",x"000026aa",x"000026ab",x"000026ab",x"000026ac",x"000026ad",x"000026ad",
		x"000026ae",x"000026af",x"000026af",x"000026b0",x"000026b0",x"000026b1",x"000026b2",x"000026b2",
		x"000026b3",x"000026b3",x"000026b4",x"000026b5",x"000026b5",x"000026b6",x"000026b6",x"000026b7",
		x"000026b8",x"000026b8",x"000026b9",x"000026b9",x"000026ba",x"000026ba",x"000026bb",x"000026bc",
		x"000026bc",x"000026bd",x"000026bd",x"000026be",x"000026be",x"000026bf",x"000026c0",x"000026c0",
		x"000026c1",x"000026c1",x"000026c2",x"000026c2",x"000026c3",x"000026c3",x"000026c4",x"000026c5",
		x"000026c5",x"000026c6",x"000026c6",x"000026c7",x"000026c7",x"000026c8",x"000026c8",x"000026c9",
		x"000026c9",x"000026ca",x"000026ca",x"000026cb",x"000026cb",x"000026cc",x"000026cd",x"000026cd",
		x"000026ce",x"000026ce",x"000026cf",x"000026cf",x"000026d0",x"000026d0",x"000026d1",x"000026d1",
		x"000026d2",x"000026d2",x"000026d3",x"000026d3",x"000026d4",x"000026d4",x"000026d5",x"000026d5",
		x"000026d5",x"000026d6",x"000026d6",x"000026d7",x"000026d7",x"000026d8",x"000026d8",x"000026d9",
		x"000026d9",x"000026da",x"000026da",x"000026db",x"000026db",x"000026dc",x"000026dc",x"000026dc",
		x"000026dd",x"000026dd",x"000026de",x"000026de",x"000026df",x"000026df",x"000026e0",x"000026e0",
		x"000026e0",x"000026e1",x"000026e1",x"000026e2",x"000026e2",x"000026e3",x"000026e3",x"000026e3",
		x"000026e4",x"000026e4",x"000026e5",x"000026e5",x"000026e5",x"000026e6",x"000026e6",x"000026e7",
		x"000026e7",x"000026e7",x"000026e8",x"000026e8",x"000026e9",x"000026e9",x"000026e9",x"000026ea",
		x"000026ea",x"000026eb",x"000026eb",x"000026eb",x"000026ec",x"000026ec",x"000026ec",x"000026ed",
		x"000026ed",x"000026ee",x"000026ee",x"000026ee",x"000026ef",x"000026ef",x"000026ef",x"000026f0",
		x"000026f0",x"000026f0",x"000026f1",x"000026f1",x"000026f2",x"000026f2",x"000026f2",x"000026f3",
		x"000026f3",x"000026f3",x"000026f4",x"000026f4",x"000026f4",x"000026f5",x"000026f5",x"000026f5",
		x"000026f6",x"000026f6",x"000026f6",x"000026f7",x"000026f7",x"000026f7",x"000026f7",x"000026f8",
		x"000026f8",x"000026f8",x"000026f9",x"000026f9",x"000026f9",x"000026fa",x"000026fa",x"000026fa",
		x"000026fa",x"000026fb",x"000026fb",x"000026fb",x"000026fc",x"000026fc",x"000026fc",x"000026fc",
		x"000026fd",x"000026fd",x"000026fd",x"000026fe",x"000026fe",x"000026fe",x"000026fe",x"000026ff",
		x"000026ff",x"000026ff",x"000026ff",x"00002700",x"00002700",x"00002700",x"00002700",x"00002701",
		x"00002701",x"00002701",x"00002701",x"00002702",x"00002702",x"00002702",x"00002702",x"00002703",
		x"00002703",x"00002703",x"00002703",x"00002703",x"00002704",x"00002704",x"00002704",x"00002704",
		x"00002705",x"00002705",x"00002705",x"00002705",x"00002705",x"00002706",x"00002706",x"00002706",
		x"00002706",x"00002706",x"00002707",x"00002707",x"00002707",x"00002707",x"00002707",x"00002708",
		x"00002708",x"00002708",x"00002708",x"00002708",x"00002708",x"00002709",x"00002709",x"00002709",
		x"00002709",x"00002709",x"00002709",x"0000270a",x"0000270a",x"0000270a",x"0000270a",x"0000270a",
		x"0000270a",x"0000270a",x"0000270b",x"0000270b",x"0000270b",x"0000270b",x"0000270b",x"0000270b",
		x"0000270b",x"0000270c",x"0000270c",x"0000270c",x"0000270c",x"0000270c",x"0000270c",x"0000270c",
		x"0000270c",x"0000270d",x"0000270d",x"0000270d",x"0000270d",x"0000270d",x"0000270d",x"0000270d",
		x"0000270d",x"0000270d",x"0000270e",x"0000270e",x"0000270e",x"0000270e",x"0000270e",x"0000270e",
		x"0000270e",x"0000270e",x"0000270e",x"0000270e",x"0000270e",x"0000270f",x"0000270f",x"0000270f",
		x"0000270f",x"0000270f",x"0000270f",x"0000270f",x"0000270f",x"0000270f",x"0000270f",x"0000270f",
		x"0000270f",x"0000270f",x"0000270f",x"0000270f",x"0000270f",x"0000270f",x"00002710",x"00002710",
		x"00002710",x"00002710",x"00002710",x"00002710",x"00002710",x"00002710",x"00002710",x"00002710",
		x"00002710",x"00002710",x"00002710",x"00002710",x"00002710",x"00002710",x"00002710",x"00002710",
		x"00002710",x"00002710",x"00002710",x"00002710",x"00002710",x"00002710",x"00002710",x"00002710",
		x"00002710",x"00002710",x"00002710",x"00002710",x"00002710",x"00002710",x"00002710",x"00002710",
		x"00002710",x"00002710",x"00002710",x"00002710",x"00002710",x"00002710",x"00002710",x"00002710",
		x"00002710",x"00002710",x"00002710",x"0000270f",x"0000270f",x"0000270f",x"0000270f",x"0000270f",
		x"0000270f",x"0000270f",x"0000270f",x"0000270f",x"0000270f",x"0000270f",x"0000270f",x"0000270f",
		x"0000270f",x"0000270f",x"0000270f",x"0000270e",x"0000270e",x"0000270e",x"0000270e",x"0000270e",
		x"0000270e",x"0000270e",x"0000270e",x"0000270e",x"0000270e",x"0000270e",x"0000270e",x"0000270d",
		x"0000270d",x"0000270d",x"0000270d",x"0000270d",x"0000270d",x"0000270d",x"0000270d",x"0000270d",
		x"0000270c",x"0000270c",x"0000270c",x"0000270c",x"0000270c",x"0000270c",x"0000270c",x"0000270c",
		x"0000270b",x"0000270b",x"0000270b",x"0000270b",x"0000270b",x"0000270b",x"0000270b",x"0000270a",
		x"0000270a",x"0000270a",x"0000270a",x"0000270a",x"0000270a",x"00002709",x"00002709",x"00002709",
		x"00002709",x"00002709",x"00002709",x"00002708",x"00002708",x"00002708",x"00002708",x"00002708",
		x"00002708",x"00002707",x"00002707",x"00002707",x"00002707",x"00002707",x"00002706",x"00002706",
		x"00002706",x"00002706",x"00002706",x"00002705",x"00002705",x"00002705",x"00002705",x"00002705",
		x"00002704",x"00002704",x"00002704",x"00002704",x"00002704",x"00002703",x"00002703",x"00002703",
		x"00002703",x"00002702",x"00002702",x"00002702",x"00002702",x"00002701",x"00002701",x"00002701",
		x"00002701",x"00002701",x"00002700",x"00002700",x"00002700",x"00002700",x"000026ff",x"000026ff",
		x"000026ff",x"000026fe",x"000026fe",x"000026fe",x"000026fe",x"000026fd",x"000026fd",x"000026fd",
		x"000026fd",x"000026fc",x"000026fc",x"000026fc",x"000026fb",x"000026fb",x"000026fb",x"000026fb",
		x"000026fa",x"000026fa",x"000026fa",x"000026f9",x"000026f9",x"000026f9",x"000026f9",x"000026f8",
		x"000026f8",x"000026f8",x"000026f7",x"000026f7",x"000026f7",x"000026f6",x"000026f6",x"000026f6",
		x"000026f5",x"000026f5",x"000026f5",x"000026f4",x"000026f4",x"000026f4",x"000026f3",x"000026f3",
		x"000026f3",x"000026f2",x"000026f2",x"000026f2",x"000026f1",x"000026f1",x"000026f1",x"000026f0",
		x"000026f0",x"000026f0",x"000026ef",x"000026ef",x"000026ef",x"000026ee",x"000026ee",x"000026ed",
		x"000026ed",x"000026ed",x"000026ec",x"000026ec",x"000026ec",x"000026eb",x"000026eb",x"000026ea",
		x"000026ea",x"000026ea",x"000026e9",x"000026e9",x"000026e8",x"000026e8",x"000026e8",x"000026e7",
		x"000026e7",x"000026e6",x"000026e6",x"000026e6",x"000026e5",x"000026e5",x"000026e4",x"000026e4",
		x"000026e4",x"000026e3",x"000026e3",x"000026e2",x"000026e2",x"000026e1",x"000026e1",x"000026e1",
		x"000026e0",x"000026e0",x"000026df",x"000026df",x"000026de",x"000026de",x"000026de",x"000026dd",
		x"000026dd",x"000026dc",x"000026dc",x"000026db",x"000026db",x"000026da",x"000026da",x"000026d9",
		x"000026d9",x"000026d9",x"000026d8",x"000026d8",x"000026d7",x"000026d7",x"000026d6",x"000026d6",
		x"000026d5",x"000026d5",x"000026d4",x"000026d4",x"000026d3",x"000026d3",x"000026d2",x"000026d2",
		x"000026d1",x"000026d1",x"000026d0",x"000026d0",x"000026cf",x"000026cf",x"000026ce",x"000026ce",
		x"000026cd",x"000026cd",x"000026cc",x"000026cc",x"000026cb",x"000026cb",x"000026ca",x"000026ca",
		x"000026c9",x"000026c9",x"000026c8",x"000026c8",x"000026c7",x"000026c6",x"000026c6",x"000026c5",
		x"000026c5",x"000026c4",x"000026c4",x"000026c3",x"000026c3",x"000026c2",x"000026c2",x"000026c1",
		x"000026c0",x"000026c0",x"000026bf",x"000026bf",x"000026be",x"000026be",x"000026bd",x"000026bc",
		x"000026bc",x"000026bb",x"000026bb",x"000026ba",x"000026ba",x"000026b9",x"000026b8",x"000026b8",
		x"000026b7",x"000026b7",x"000026b6",x"000026b5",x"000026b5",x"000026b4",x"000026b4",x"000026b3",
		x"000026b2",x"000026b2",x"000026b1",x"000026b1",x"000026b0",x"000026af",x"000026af",x"000026ae",
		x"000026ae",x"000026ad",x"000026ac",x"000026ac",x"000026ab",x"000026aa",x"000026aa",x"000026a9",
		x"000026a9",x"000026a8",x"000026a7",x"000026a7",x"000026a6",x"000026a5",x"000026a5",x"000026a4",
		x"000026a3",x"000026a3",x"000026a2",x"000026a1",x"000026a1",x"000026a0",x"0000269f",x"0000269f",
		x"0000269e",x"0000269d",x"0000269d",x"0000269c",x"0000269b",x"0000269b",x"0000269a",x"00002699",
		x"00002699",x"00002698",x"00002697",x"00002697",x"00002696",x"00002695",x"00002695",x"00002694",
		x"00002693",x"00002693",x"00002692",x"00002691",x"00002690",x"00002690",x"0000268f",x"0000268e",
		x"0000268e",x"0000268d",x"0000268c",x"0000268b",x"0000268b",x"0000268a",x"00002689",x"00002689",
		x"00002688",x"00002687",x"00002686",x"00002686",x"00002685",x"00002684",x"00002683",x"00002683",
		x"00002682",x"00002681",x"00002680",x"00002680",x"0000267f",x"0000267e",x"0000267d",x"0000267d",
		x"0000267c",x"0000267b",x"0000267a",x"0000267a",x"00002679",x"00002678",x"00002677",x"00002677",
		x"00002676",x"00002675",x"00002674",x"00002673",x"00002673",x"00002672",x"00002671",x"00002670",
		x"00002670",x"0000266f",x"0000266e",x"0000266d",x"0000266c",x"0000266c",x"0000266b",x"0000266a",
		x"00002669",x"00002668",x"00002668",x"00002667",x"00002666",x"00002665",x"00002664",x"00002663",
		x"00002663",x"00002662",x"00002661",x"00002660",x"0000265f",x"0000265f",x"0000265e",x"0000265d",
		x"0000265c",x"0000265b",x"0000265a",x"0000265a",x"00002659",x"00002658",x"00002657",x"00002656",
		x"00002655",x"00002654",x"00002654",x"00002653",x"00002652",x"00002651",x"00002650",x"0000264f",
		x"0000264e",x"0000264e",x"0000264d",x"0000264c",x"0000264b",x"0000264a",x"00002649",x"00002648",
		x"00002647",x"00002647",x"00002646",x"00002645",x"00002644",x"00002643",x"00002642",x"00002641",
		x"00002640",x"0000263f",x"0000263f",x"0000263e",x"0000263d",x"0000263c",x"0000263b",x"0000263a",
		x"00002639",x"00002638",x"00002637",x"00002636",x"00002635",x"00002635",x"00002634",x"00002633",
		x"00002632",x"00002631",x"00002630",x"0000262f",x"0000262e",x"0000262d",x"0000262c",x"0000262b",
		x"0000262a",x"00002629",x"00002628",x"00002627",x"00002627",x"00002626",x"00002625",x"00002624",
		x"00002623",x"00002622",x"00002621",x"00002620",x"0000261f",x"0000261e",x"0000261d",x"0000261c",
		x"0000261b",x"0000261a",x"00002619",x"00002618",x"00002617",x"00002616",x"00002615",x"00002614",
		x"00002613",x"00002612",x"00002611",x"00002610",x"0000260f",x"0000260e",x"0000260d",x"0000260c",
		x"0000260b",x"0000260a",x"00002609",x"00002608",x"00002607",x"00002606",x"00002605",x"00002604",
		x"00002603",x"00002602",x"00002601",x"00002600",x"000025ff",x"000025fe",x"000025fd",x"000025fc",
		x"000025fb",x"000025fa",x"000025f9",x"000025f8",x"000025f7",x"000025f6",x"000025f5",x"000025f4",
		x"000025f3",x"000025f2",x"000025f1",x"000025ef",x"000025ee",x"000025ed",x"000025ec",x"000025eb",
		x"000025ea",x"000025e9",x"000025e8",x"000025e7",x"000025e6",x"000025e5",x"000025e4",x"000025e3",
		x"000025e2",x"000025e1",x"000025e0",x"000025de",x"000025dd",x"000025dc",x"000025db",x"000025da",
		x"000025d9",x"000025d8",x"000025d7",x"000025d6",x"000025d5",x"000025d4",x"000025d2",x"000025d1",
		x"000025d0",x"000025cf",x"000025ce",x"000025cd",x"000025cc",x"000025cb",x"000025ca",x"000025c8",
		x"000025c7",x"000025c6",x"000025c5",x"000025c4",x"000025c3",x"000025c2",x"000025c1",x"000025bf",
		x"000025be",x"000025bd",x"000025bc",x"000025bb",x"000025ba",x"000025b9",x"000025b7",x"000025b6",
		x"000025b5",x"000025b4",x"000025b3",x"000025b2",x"000025b1",x"000025af",x"000025ae",x"000025ad",
		x"000025ac",x"000025ab",x"000025aa",x"000025a8",x"000025a7",x"000025a6",x"000025a5",x"000025a4",
		x"000025a3",x"000025a1",x"000025a0",x"0000259f",x"0000259e",x"0000259d",x"0000259b",x"0000259a",
		x"00002599",x"00002598",x"00002597",x"00002595",x"00002594",x"00002593",x"00002592",x"00002591",
		x"0000258f",x"0000258e",x"0000258d",x"0000258c",x"0000258b",x"00002589",x"00002588",x"00002587",
		x"00002586",x"00002584",x"00002583",x"00002582",x"00002581",x"00002580",x"0000257e",x"0000257d",
		x"0000257c",x"0000257b",x"00002579",x"00002578",x"00002577",x"00002576",x"00002574",x"00002573",
		x"00002572",x"00002571",x"0000256f",x"0000256e",x"0000256d",x"0000256c",x"0000256a",x"00002569",
		x"00002568",x"00002567",x"00002565",x"00002564",x"00002563",x"00002561",x"00002560",x"0000255f",
		x"0000255e",x"0000255c",x"0000255b",x"0000255a",x"00002558",x"00002557",x"00002556",x"00002555",
		x"00002553",x"00002552",x"00002551",x"0000254f",x"0000254e",x"0000254d",x"0000254c",x"0000254a",
		x"00002549",x"00002548",x"00002546",x"00002545",x"00002544",x"00002542",x"00002541",x"00002540",
		x"0000253e",x"0000253d",x"0000253c",x"0000253a",x"00002539",x"00002538",x"00002536",x"00002535",
		x"00002534",x"00002532",x"00002531",x"00002530",x"0000252e",x"0000252d",x"0000252c",x"0000252a",
		x"00002529",x"00002528",x"00002526",x"00002525",x"00002524",x"00002522",x"00002521",x"0000251f",
		x"0000251e",x"0000251d",x"0000251b",x"0000251a",x"00002519",x"00002517",x"00002516",x"00002514",
		x"00002513",x"00002512",x"00002510",x"0000250f",x"0000250e",x"0000250c",x"0000250b",x"00002509",
		x"00002508",x"00002507",x"00002505",x"00002504",x"00002502",x"00002501",x"00002500",x"000024fe",
		x"000024fd",x"000024fb",x"000024fa",x"000024f9",x"000024f7",x"000024f6",x"000024f4",x"000024f3",
		x"000024f1",x"000024f0",x"000024ef",x"000024ed",x"000024ec",x"000024ea",x"000024e9",x"000024e7",
		x"000024e6",x"000024e5",x"000024e3",x"000024e2",x"000024e0",x"000024df",x"000024dd",x"000024dc",
		x"000024da",x"000024d9",x"000024d8",x"000024d6",x"000024d5",x"000024d3",x"000024d2",x"000024d0",
		x"000024cf",x"000024cd",x"000024cc",x"000024ca",x"000024c9",x"000024c7",x"000024c6",x"000024c4",
		x"000024c3",x"000024c1",x"000024c0",x"000024bf",x"000024bd",x"000024bc",x"000024ba",x"000024b9",
		x"000024b7",x"000024b6",x"000024b4",x"000024b3",x"000024b1",x"000024b0",x"000024ae",x"000024ad",
		x"000024ab",x"000024aa",x"000024a8",x"000024a7",x"000024a5",x"000024a4",x"000024a2",x"000024a0",
		x"0000249f",x"0000249d",x"0000249c",x"0000249a",x"00002499",x"00002497",x"00002496",x"00002494",
		x"00002493",x"00002491",x"00002490",x"0000248e",x"0000248d",x"0000248b",x"00002489",x"00002488",
		x"00002486",x"00002485",x"00002483",x"00002482",x"00002480",x"0000247f",x"0000247d",x"0000247c",
		x"0000247a",x"00002478",x"00002477",x"00002475",x"00002474",x"00002472",x"00002471",x"0000246f",
		x"0000246d",x"0000246c",x"0000246a",x"00002469",x"00002467",x"00002466",x"00002464",x"00002462",
		x"00002461",x"0000245f",x"0000245e",x"0000245c",x"0000245a",x"00002459",x"00002457",x"00002456",
		x"00002454",x"00002452",x"00002451",x"0000244f",x"0000244e",x"0000244c",x"0000244a",x"00002449",
		x"00002447",x"00002445",x"00002444",x"00002442",x"00002441",x"0000243f",x"0000243d",x"0000243c",
		x"0000243a",x"00002438",x"00002437",x"00002435",x"00002434",x"00002432",x"00002430",x"0000242f",
		x"0000242d",x"0000242b",x"0000242a",x"00002428",x"00002426",x"00002425",x"00002423",x"00002421",
		x"00002420",x"0000241e",x"0000241c",x"0000241b",x"00002419",x"00002417",x"00002416",x"00002414",
		x"00002412",x"00002411",x"0000240f",x"0000240d",x"0000240c",x"0000240a",x"00002408",x"00002407",
		x"00002405",x"00002403",x"00002402",x"00002400",x"000023fe",x"000023fd",x"000023fb",x"000023f9",
		x"000023f8",x"000023f6",x"000023f4",x"000023f2",x"000023f1",x"000023ef",x"000023ed",x"000023ec",
		x"000023ea",x"000023e8",x"000023e6",x"000023e5",x"000023e3",x"000023e1",x"000023e0",x"000023de",
		x"000023dc",x"000023da",x"000023d9",x"000023d7",x"000023d5",x"000023d4",x"000023d2",x"000023d0",
		x"000023ce",x"000023cd",x"000023cb",x"000023c9",x"000023c7",x"000023c6",x"000023c4",x"000023c2",
		x"000023c0",x"000023bf",x"000023bd",x"000023bb",x"000023b9",x"000023b8",x"000023b6",x"000023b4",
		x"000023b2",x"000023b1",x"000023af",x"000023ad",x"000023ab",x"000023a9",x"000023a8",x"000023a6",
		x"000023a4",x"000023a2",x"000023a1",x"0000239f",x"0000239d",x"0000239b",x"00002399",x"00002398",
		x"00002396",x"00002394",x"00002392",x"00002391",x"0000238f",x"0000238d",x"0000238b",x"00002389",
		x"00002388",x"00002386",x"00002384",x"00002382",x"00002380",x"0000237f",x"0000237d",x"0000237b",
		x"00002379",x"00002377",x"00002375",x"00002374",x"00002372",x"00002370",x"0000236e",x"0000236c",
		x"0000236a",x"00002369",x"00002367",x"00002365",x"00002363",x"00002361",x"0000235f",x"0000235e",
		x"0000235c",x"0000235a",x"00002358",x"00002356",x"00002354",x"00002353",x"00002351",x"0000234f",
		x"0000234d",x"0000234b",x"00002349",x"00002347",x"00002346",x"00002344",x"00002342",x"00002340",
		x"0000233e",x"0000233c",x"0000233a",x"00002339",x"00002337",x"00002335",x"00002333",x"00002331",
		x"0000232f",x"0000232d",x"0000232b",x"0000232a",x"00002328",x"00002326",x"00002324",x"00002322",
		x"00002320",x"0000231e",x"0000231c",x"0000231a",x"00002319",x"00002317",x"00002315",x"00002313",
		x"00002311",x"0000230f",x"0000230d",x"0000230b",x"00002309",x"00002307",x"00002305",x"00002304",
		x"00002302",x"00002300",x"000022fe",x"000022fc",x"000022fa",x"000022f8",x"000022f6",x"000022f4",
		x"000022f2",x"000022f0",x"000022ee",x"000022ec",x"000022eb",x"000022e9",x"000022e7",x"000022e5",
		x"000022e3",x"000022e1",x"000022df",x"000022dd",x"000022db",x"000022d9",x"000022d7",x"000022d5",
		x"000022d3",x"000022d1",x"000022cf",x"000022cd",x"000022cb",x"000022c9",x"000022c7",x"000022c5",
		x"000022c3",x"000022c2",x"000022c0",x"000022be",x"000022bc",x"000022ba",x"000022b8",x"000022b6",
		x"000022b4",x"000022b2",x"000022b0",x"000022ae",x"000022ac",x"000022aa",x"000022a8",x"000022a6",
		x"000022a4",x"000022a2",x"000022a0",x"0000229e",x"0000229c",x"0000229a",x"00002298",x"00002296",
		x"00002294",x"00002292",x"00002290",x"0000228e",x"0000228c",x"0000228a",x"00002288",x"00002286",
		x"00002284",x"00002282",x"00002280",x"0000227e",x"0000227c",x"0000227a",x"00002278",x"00002276",
		x"00002274",x"00002272",x"00002270",x"0000226e",x"0000226b",x"00002269",x"00002267",x"00002265",
		x"00002263",x"00002261",x"0000225f",x"0000225d",x"0000225b",x"00002259",x"00002257",x"00002255",
		x"00002253",x"00002251",x"0000224f",x"0000224d",x"0000224b",x"00002249",x"00002247",x"00002245",
		x"00002243",x"00002240",x"0000223e",x"0000223c",x"0000223a",x"00002238",x"00002236",x"00002234",
		x"00002232",x"00002230",x"0000222e",x"0000222c",x"0000222a",x"00002228",x"00002225",x"00002223",
		x"00002221",x"0000221f",x"0000221d",x"0000221b",x"00002219",x"00002217",x"00002215",x"00002213",
		x"00002211",x"0000220e",x"0000220c",x"0000220a",x"00002208",x"00002206",x"00002204",x"00002202",
		x"00002200",x"000021fe",x"000021fb",x"000021f9",x"000021f7",x"000021f5",x"000021f3",x"000021f1",
		x"000021ef",x"000021ed",x"000021eb",x"000021e8",x"000021e6",x"000021e4",x"000021e2",x"000021e0",
		x"000021de",x"000021dc",x"000021d9",x"000021d7",x"000021d5",x"000021d3",x"000021d1",x"000021cf",
		x"000021cd",x"000021ca",x"000021c8",x"000021c6",x"000021c4",x"000021c2",x"000021c0",x"000021be",
		x"000021bb",x"000021b9",x"000021b7",x"000021b5",x"000021b3",x"000021b1",x"000021ae",x"000021ac",
		x"000021aa",x"000021a8",x"000021a6",x"000021a4",x"000021a1",x"0000219f",x"0000219d",x"0000219b",
		x"00002199",x"00002197",x"00002194",x"00002192",x"00002190",x"0000218e",x"0000218c",x"00002189",
		x"00002187",x"00002185",x"00002183",x"00002181",x"0000217e",x"0000217c",x"0000217a",x"00002178",
		x"00002176",x"00002173",x"00002171",x"0000216f",x"0000216d",x"0000216b",x"00002168",x"00002166",
		x"00002164",x"00002162",x"00002160",x"0000215d",x"0000215b",x"00002159",x"00002157",x"00002154",
		x"00002152",x"00002150",x"0000214e",x"0000214c",x"00002149",x"00002147",x"00002145",x"00002143",
		x"00002140",x"0000213e",x"0000213c",x"0000213a",x"00002137",x"00002135",x"00002133",x"00002131",
		x"0000212e",x"0000212c",x"0000212a",x"00002128",x"00002125",x"00002123",x"00002121",x"0000211f",
		x"0000211c",x"0000211a",x"00002118",x"00002116",x"00002113",x"00002111",x"0000210f",x"0000210d",
		x"0000210a",x"00002108",x"00002106",x"00002104",x"00002101",x"000020ff",x"000020fd",x"000020fa",
		x"000020f8",x"000020f6",x"000020f4",x"000020f1",x"000020ef",x"000020ed",x"000020ea",x"000020e8",
		x"000020e6",x"000020e4",x"000020e1",x"000020df",x"000020dd",x"000020da",x"000020d8",x"000020d6",
		x"000020d3",x"000020d1",x"000020cf",x"000020cd",x"000020ca",x"000020c8",x"000020c6",x"000020c3",
		x"000020c1",x"000020bf",x"000020bc",x"000020ba",x"000020b8",x"000020b5",x"000020b3",x"000020b1",
		x"000020ae",x"000020ac",x"000020aa",x"000020a8",x"000020a5",x"000020a3",x"000020a1",x"0000209e",
		x"0000209c",x"0000209a",x"00002097",x"00002095",x"00002093",x"00002090",x"0000208e",x"0000208c",
		x"00002089",x"00002087",x"00002084",x"00002082",x"00002080",x"0000207d",x"0000207b",x"00002079",
		x"00002076",x"00002074",x"00002072",x"0000206f",x"0000206d",x"0000206b",x"00002068",x"00002066",
		x"00002063",x"00002061",x"0000205f",x"0000205c",x"0000205a",x"00002058",x"00002055",x"00002053",
		x"00002051",x"0000204e",x"0000204c",x"00002049",x"00002047",x"00002045",x"00002042",x"00002040",
		x"0000203d",x"0000203b",x"00002039",x"00002036",x"00002034",x"00002032",x"0000202f",x"0000202d",
		x"0000202a",x"00002028",x"00002026",x"00002023",x"00002021",x"0000201e",x"0000201c",x"0000201a",
		x"00002017",x"00002015",x"00002012",x"00002010",x"0000200e",x"0000200b",x"00002009",x"00002006",
		x"00002004",x"00002001",x"00001fff",x"00001ffd",x"00001ffa",x"00001ff8",x"00001ff5",x"00001ff3",
		x"00001ff0",x"00001fee",x"00001fec",x"00001fe9",x"00001fe7",x"00001fe4",x"00001fe2",x"00001fdf",
		x"00001fdd",x"00001fdb",x"00001fd8",x"00001fd6",x"00001fd3",x"00001fd1",x"00001fce",x"00001fcc",
		x"00001fc9",x"00001fc7",x"00001fc5",x"00001fc2",x"00001fc0",x"00001fbd",x"00001fbb",x"00001fb8",
		x"00001fb6",x"00001fb3",x"00001fb1",x"00001faf",x"00001fac",x"00001faa",x"00001fa7",x"00001fa5",
		x"00001fa2",x"00001fa0",x"00001f9d",x"00001f9b",x"00001f98",x"00001f96",x"00001f93",x"00001f91",
		x"00001f8e",x"00001f8c",x"00001f89",x"00001f87",x"00001f85",x"00001f82",x"00001f80",x"00001f7d",
		x"00001f7b",x"00001f78",x"00001f76",x"00001f73",x"00001f71",x"00001f6e",x"00001f6c",x"00001f69",
		x"00001f67",x"00001f64",x"00001f62",x"00001f5f",x"00001f5d",x"00001f5a",x"00001f58",x"00001f55",
		x"00001f53",x"00001f50",x"00001f4e",x"00001f4b",x"00001f49",x"00001f46",x"00001f44",x"00001f41",
		x"00001f3f",x"00001f3c",x"00001f3a",x"00001f37",x"00001f35",x"00001f32",x"00001f2f",x"00001f2d",
		x"00001f2a",x"00001f28",x"00001f25",x"00001f23",x"00001f20",x"00001f1e",x"00001f1b",x"00001f19",
		x"00001f16",x"00001f14",x"00001f11",x"00001f0f",x"00001f0c",x"00001f0a",x"00001f07",x"00001f04",
		x"00001f02",x"00001eff",x"00001efd",x"00001efa",x"00001ef8",x"00001ef5",x"00001ef3",x"00001ef0",
		x"00001eee",x"00001eeb",x"00001ee8",x"00001ee6",x"00001ee3",x"00001ee1",x"00001ede",x"00001edc",
		x"00001ed9",x"00001ed7",x"00001ed4",x"00001ed1",x"00001ecf",x"00001ecc",x"00001eca",x"00001ec7",
		x"00001ec5",x"00001ec2",x"00001ebf",x"00001ebd",x"00001eba",x"00001eb8",x"00001eb5",x"00001eb3",
		x"00001eb0",x"00001ead",x"00001eab",x"00001ea8",x"00001ea6",x"00001ea3",x"00001ea0",x"00001e9e",
		x"00001e9b",x"00001e99",x"00001e96",x"00001e94",x"00001e91",x"00001e8e",x"00001e8c",x"00001e89",
		x"00001e87",x"00001e84",x"00001e81",x"00001e7f",x"00001e7c",x"00001e7a",x"00001e77",x"00001e74",
		x"00001e72",x"00001e6f",x"00001e6d",x"00001e6a",x"00001e67",x"00001e65",x"00001e62",x"00001e5f",
		x"00001e5d",x"00001e5a",x"00001e58",x"00001e55",x"00001e52",x"00001e50",x"00001e4d",x"00001e4b",
		x"00001e48",x"00001e45",x"00001e43",x"00001e40",x"00001e3d",x"00001e3b",x"00001e38",x"00001e36",
		x"00001e33",x"00001e30",x"00001e2e",x"00001e2b",x"00001e28",x"00001e26",x"00001e23",x"00001e20",
		x"00001e1e",x"00001e1b",x"00001e19",x"00001e16",x"00001e13",x"00001e11",x"00001e0e",x"00001e0b",
		x"00001e09",x"00001e06",x"00001e03",x"00001e01",x"00001dfe",x"00001dfb",x"00001df9",x"00001df6",
		x"00001df3",x"00001df1",x"00001dee",x"00001deb",x"00001de9",x"00001de6",x"00001de3",x"00001de1",
		x"00001dde",x"00001ddb",x"00001dd9",x"00001dd6",x"00001dd3",x"00001dd1",x"00001dce",x"00001dcb",
		x"00001dc9",x"00001dc6",x"00001dc3",x"00001dc1",x"00001dbe",x"00001dbb",x"00001db9",x"00001db6",
		x"00001db3",x"00001db1",x"00001dae",x"00001dab",x"00001da9",x"00001da6",x"00001da3",x"00001da1",
		x"00001d9e",x"00001d9b",x"00001d98",x"00001d96",x"00001d93",x"00001d90",x"00001d8e",x"00001d8b",
		x"00001d88",x"00001d86",x"00001d83",x"00001d80",x"00001d7d",x"00001d7b",x"00001d78",x"00001d75",
		x"00001d73",x"00001d70",x"00001d6d",x"00001d6b",x"00001d68",x"00001d65",x"00001d62",x"00001d60",
		x"00001d5d",x"00001d5a",x"00001d58",x"00001d55",x"00001d52",x"00001d4f",x"00001d4d",x"00001d4a",
		x"00001d47",x"00001d45",x"00001d42",x"00001d3f",x"00001d3c",x"00001d3a",x"00001d37",x"00001d34",
		x"00001d31",x"00001d2f",x"00001d2c",x"00001d29",x"00001d26",x"00001d24",x"00001d21",x"00001d1e",
		x"00001d1c",x"00001d19",x"00001d16",x"00001d13",x"00001d11",x"00001d0e",x"00001d0b",x"00001d08",
		x"00001d06",x"00001d03",x"00001d00",x"00001cfd",x"00001cfb",x"00001cf8",x"00001cf5",x"00001cf2",
		x"00001cf0",x"00001ced",x"00001cea",x"00001ce7",x"00001ce5",x"00001ce2",x"00001cdf",x"00001cdc",
		x"00001cda",x"00001cd7",x"00001cd4",x"00001cd1",x"00001cce",x"00001ccc",x"00001cc9",x"00001cc6",
		x"00001cc3",x"00001cc1",x"00001cbe",x"00001cbb",x"00001cb8",x"00001cb6",x"00001cb3",x"00001cb0",
		x"00001cad",x"00001caa",x"00001ca8",x"00001ca5",x"00001ca2",x"00001c9f",x"00001c9d",x"00001c9a",
		x"00001c97",x"00001c94",x"00001c91",x"00001c8f",x"00001c8c",x"00001c89",x"00001c86",x"00001c84",
		x"00001c81",x"00001c7e",x"00001c7b",x"00001c78",x"00001c76",x"00001c73",x"00001c70",x"00001c6d",
		x"00001c6a",x"00001c68",x"00001c65",x"00001c62",x"00001c5f",x"00001c5c",x"00001c5a",x"00001c57",
		x"00001c54",x"00001c51",x"00001c4e",x"00001c4c",x"00001c49",x"00001c46",x"00001c43",x"00001c40",
		x"00001c3d",x"00001c3b",x"00001c38",x"00001c35",x"00001c32",x"00001c2f",x"00001c2d",x"00001c2a",
		x"00001c27",x"00001c24",x"00001c21",x"00001c1e",x"00001c1c",x"00001c19",x"00001c16",x"00001c13",
		x"00001c10",x"00001c0e",x"00001c0b",x"00001c08",x"00001c05",x"00001c02",x"00001bff",x"00001bfd",
		x"00001bfa",x"00001bf7",x"00001bf4",x"00001bf1",x"00001bee",x"00001bec",x"00001be9",x"00001be6",
		x"00001be3",x"00001be0",x"00001bdd",x"00001bdb",x"00001bd8",x"00001bd5",x"00001bd2",x"00001bcf",
		x"00001bcc",x"00001bc9",x"00001bc7",x"00001bc4",x"00001bc1",x"00001bbe",x"00001bbb",x"00001bb8",
		x"00001bb5",x"00001bb3",x"00001bb0",x"00001bad",x"00001baa",x"00001ba7",x"00001ba4",x"00001ba2",
		x"00001b9f",x"00001b9c",x"00001b99",x"00001b96",x"00001b93",x"00001b90",x"00001b8d",x"00001b8b",
		x"00001b88",x"00001b85",x"00001b82",x"00001b7f",x"00001b7c",x"00001b79",x"00001b77",x"00001b74",
		x"00001b71",x"00001b6e",x"00001b6b",x"00001b68",x"00001b65",x"00001b62",x"00001b60",x"00001b5d",
		x"00001b5a",x"00001b57",x"00001b54",x"00001b51",x"00001b4e",x"00001b4b",x"00001b48",x"00001b46",
		x"00001b43",x"00001b40",x"00001b3d",x"00001b3a",x"00001b37",x"00001b34",x"00001b31",x"00001b2e",
		x"00001b2c",x"00001b29",x"00001b26",x"00001b23",x"00001b20",x"00001b1d",x"00001b1a",x"00001b17",
		x"00001b14",x"00001b12",x"00001b0f",x"00001b0c",x"00001b09",x"00001b06",x"00001b03",x"00001b00",
		x"00001afd",x"00001afa",x"00001af7",x"00001af5",x"00001af2",x"00001aef",x"00001aec",x"00001ae9",
		x"00001ae6",x"00001ae3",x"00001ae0",x"00001add",x"00001ada",x"00001ad7",x"00001ad5",x"00001ad2",
		x"00001acf",x"00001acc",x"00001ac9",x"00001ac6",x"00001ac3",x"00001ac0",x"00001abd",x"00001aba",
		x"00001ab7",x"00001ab4",x"00001ab1",x"00001aaf",x"00001aac",x"00001aa9",x"00001aa6",x"00001aa3",
		x"00001aa0",x"00001a9d",x"00001a9a",x"00001a97",x"00001a94",x"00001a91",x"00001a8e",x"00001a8b",
		x"00001a88",x"00001a86",x"00001a83",x"00001a80",x"00001a7d",x"00001a7a",x"00001a77",x"00001a74",
		x"00001a71",x"00001a6e",x"00001a6b",x"00001a68",x"00001a65",x"00001a62",x"00001a5f",x"00001a5c",
		x"00001a59",x"00001a57",x"00001a54",x"00001a51",x"00001a4e",x"00001a4b",x"00001a48",x"00001a45",
		x"00001a42",x"00001a3f",x"00001a3c",x"00001a39",x"00001a36",x"00001a33",x"00001a30",x"00001a2d",
		x"00001a2a",x"00001a27",x"00001a24",x"00001a21",x"00001a1e",x"00001a1c",x"00001a19",x"00001a16",
		x"00001a13",x"00001a10",x"00001a0d",x"00001a0a",x"00001a07",x"00001a04",x"00001a01",x"000019fe",
		x"000019fb",x"000019f8",x"000019f5",x"000019f2",x"000019ef",x"000019ec",x"000019e9",x"000019e6",
		x"000019e3",x"000019e0",x"000019dd",x"000019da",x"000019d7",x"000019d4",x"000019d1",x"000019ce",
		x"000019cb",x"000019c8",x"000019c5",x"000019c2",x"000019bf",x"000019bc",x"000019ba",x"000019b7",
		x"000019b4",x"000019b1",x"000019ae",x"000019ab",x"000019a8",x"000019a5",x"000019a2",x"0000199f",
		x"0000199c",x"00001999",x"00001996",x"00001993",x"00001990",x"0000198d",x"0000198a",x"00001987",
		x"00001984",x"00001981",x"0000197e",x"0000197b",x"00001978",x"00001975",x"00001972",x"0000196f",
		x"0000196c",x"00001969",x"00001966",x"00001963",x"00001960",x"0000195d",x"0000195a",x"00001957",
		x"00001954",x"00001951",x"0000194e",x"0000194b",x"00001948",x"00001945",x"00001942",x"0000193f",
		x"0000193c",x"00001939",x"00001936",x"00001933",x"00001930",x"0000192d",x"0000192a",x"00001927",
		x"00001924",x"00001921",x"0000191e",x"0000191b",x"00001918",x"00001915",x"00001912",x"0000190f",
		x"0000190c",x"00001909",x"00001906",x"00001903",x"00001900",x"000018fd",x"000018fa",x"000018f7",
		x"000018f4",x"000018f1",x"000018ee",x"000018ea",x"000018e7",x"000018e4",x"000018e1",x"000018de",
		x"000018db",x"000018d8",x"000018d5",x"000018d2",x"000018cf",x"000018cc",x"000018c9",x"000018c6",
		x"000018c3",x"000018c0",x"000018bd",x"000018ba",x"000018b7",x"000018b4",x"000018b1",x"000018ae",
		x"000018ab",x"000018a8",x"000018a5",x"000018a2",x"0000189f",x"0000189c",x"00001899",x"00001896",
		x"00001893",x"00001890",x"0000188d",x"0000188a",x"00001887",x"00001883",x"00001880",x"0000187d",
		x"0000187a",x"00001877",x"00001874",x"00001871",x"0000186e",x"0000186b",x"00001868",x"00001865",
		x"00001862",x"0000185f",x"0000185c",x"00001859",x"00001856",x"00001853",x"00001850",x"0000184d",
		x"0000184a",x"00001847",x"00001844",x"00001841",x"0000183d",x"0000183a",x"00001837",x"00001834",
		x"00001831",x"0000182e",x"0000182b",x"00001828",x"00001825",x"00001822",x"0000181f",x"0000181c",
		x"00001819",x"00001816",x"00001813",x"00001810",x"0000180d",x"0000180a",x"00001807",x"00001803",
		x"00001800",x"000017fd",x"000017fa",x"000017f7",x"000017f4",x"000017f1",x"000017ee",x"000017eb",
		x"000017e8",x"000017e5",x"000017e2",x"000017df",x"000017dc",x"000017d9",x"000017d6",x"000017d2",
		x"000017cf",x"000017cc",x"000017c9",x"000017c6",x"000017c3",x"000017c0",x"000017bd",x"000017ba",
		x"000017b7",x"000017b4",x"000017b1",x"000017ae",x"000017ab",x"000017a8",x"000017a4",x"000017a1",
		x"0000179e",x"0000179b",x"00001798",x"00001795",x"00001792",x"0000178f",x"0000178c",x"00001789",
		x"00001786",x"00001783",x"00001780",x"0000177c",x"00001779",x"00001776",x"00001773",x"00001770",
		x"0000176d",x"0000176a",x"00001767",x"00001764",x"00001761",x"0000175e",x"0000175b",x"00001758",
		x"00001754",x"00001751",x"0000174e",x"0000174b",x"00001748",x"00001745",x"00001742",x"0000173f",
		x"0000173c",x"00001739",x"00001736",x"00001733",x"0000172f",x"0000172c",x"00001729",x"00001726",
		x"00001723",x"00001720",x"0000171d",x"0000171a",x"00001717",x"00001714",x"00001711",x"0000170d",
		x"0000170a",x"00001707",x"00001704",x"00001701",x"000016fe",x"000016fb",x"000016f8",x"000016f5",
		x"000016f2",x"000016ef",x"000016eb",x"000016e8",x"000016e5",x"000016e2",x"000016df",x"000016dc",
		x"000016d9",x"000016d6",x"000016d3",x"000016d0",x"000016cd",x"000016c9",x"000016c6",x"000016c3",
		x"000016c0",x"000016bd",x"000016ba",x"000016b7",x"000016b4",x"000016b1",x"000016ae",x"000016aa",
		x"000016a7",x"000016a4",x"000016a1",x"0000169e",x"0000169b",x"00001698",x"00001695",x"00001692",
		x"0000168e",x"0000168b",x"00001688",x"00001685",x"00001682",x"0000167f",x"0000167c",x"00001679",
		x"00001676",x"00001673",x"0000166f",x"0000166c",x"00001669",x"00001666",x"00001663",x"00001660",
		x"0000165d",x"0000165a",x"00001657",x"00001653",x"00001650",x"0000164d",x"0000164a",x"00001647",
		x"00001644",x"00001641",x"0000163e",x"0000163b",x"00001637",x"00001634",x"00001631",x"0000162e",
		x"0000162b",x"00001628",x"00001625",x"00001622",x"0000161f",x"0000161b",x"00001618",x"00001615",
		x"00001612",x"0000160f",x"0000160c",x"00001609",x"00001606",x"00001603",x"000015ff",x"000015fc",
		x"000015f9",x"000015f6",x"000015f3",x"000015f0",x"000015ed",x"000015ea",x"000015e6",x"000015e3",
		x"000015e0",x"000015dd",x"000015da",x"000015d7",x"000015d4",x"000015d1",x"000015ce",x"000015ca",
		x"000015c7",x"000015c4",x"000015c1",x"000015be",x"000015bb",x"000015b8",x"000015b5",x"000015b1",
		x"000015ae",x"000015ab",x"000015a8",x"000015a5",x"000015a2",x"0000159f",x"0000159c",x"00001598",
		x"00001595",x"00001592",x"0000158f",x"0000158c",x"00001589",x"00001586",x"00001583",x"0000157f",
		x"0000157c",x"00001579",x"00001576",x"00001573",x"00001570",x"0000156d",x"0000156a",x"00001566",
		x"00001563",x"00001560",x"0000155d",x"0000155a",x"00001557",x"00001554",x"00001551",x"0000154d",
		x"0000154a",x"00001547",x"00001544",x"00001541",x"0000153e",x"0000153b",x"00001537",x"00001534",
		x"00001531",x"0000152e",x"0000152b",x"00001528",x"00001525",x"00001522",x"0000151e",x"0000151b",
		x"00001518",x"00001515",x"00001512",x"0000150f",x"0000150c",x"00001509",x"00001505",x"00001502",
		x"000014ff",x"000014fc",x"000014f9",x"000014f6",x"000014f3",x"000014ef",x"000014ec",x"000014e9",
		x"000014e6",x"000014e3",x"000014e0",x"000014dd",x"000014d9",x"000014d6",x"000014d3",x"000014d0",
		x"000014cd",x"000014ca",x"000014c7",x"000014c4",x"000014c0",x"000014bd",x"000014ba",x"000014b7",
		x"000014b4",x"000014b1",x"000014ae",x"000014aa",x"000014a7",x"000014a4",x"000014a1",x"0000149e",
		x"0000149b",x"00001498",x"00001495",x"00001491",x"0000148e",x"0000148b",x"00001488",x"00001485",
		x"00001482",x"0000147f",x"0000147b",x"00001478",x"00001475",x"00001472",x"0000146f",x"0000146c",
		x"00001469",x"00001465",x"00001462",x"0000145f",x"0000145c",x"00001459",x"00001456",x"00001453",
		x"0000144f",x"0000144c",x"00001449",x"00001446",x"00001443",x"00001440",x"0000143d",x"00001439",
		x"00001436",x"00001433",x"00001430",x"0000142d",x"0000142a",x"00001427",x"00001423",x"00001420",
		x"0000141d",x"0000141a",x"00001417",x"00001414",x"00001411",x"0000140e",x"0000140a",x"00001407",
		x"00001404",x"00001401",x"000013fe",x"000013fb",x"000013f8",x"000013f4",x"000013f1",x"000013ee",
		x"000013eb",x"000013e8",x"000013e5",x"000013e2",x"000013de",x"000013db",x"000013d8",x"000013d5",
		x"000013d2",x"000013cf",x"000013cc",x"000013c8",x"000013c5",x"000013c2",x"000013bf",x"000013bc",
		x"000013b9",x"000013b6",x"000013b2",x"000013af",x"000013ac",x"000013a9",x"000013a6",x"000013a3",
		x"000013a0",x"0000139c",x"00001399",x"00001396",x"00001393",x"00001390",x"0000138d",x"0000138a",
		x"00001386",x"00001383",x"00001380",x"0000137d",x"0000137a",x"00001377",x"00001374",x"00001370",
		x"0000136d",x"0000136a",x"00001367",x"00001364",x"00001361",x"0000135e",x"0000135a",x"00001357",
		x"00001354",x"00001351",x"0000134e",x"0000134b",x"00001348",x"00001344",x"00001341",x"0000133e",
		x"0000133b",x"00001338",x"00001335",x"00001332",x"0000132e",x"0000132b",x"00001328",x"00001325",
		x"00001322",x"0000131f",x"0000131c",x"00001318",x"00001315",x"00001312",x"0000130f",x"0000130c",
		x"00001309",x"00001306",x"00001302",x"000012ff",x"000012fc",x"000012f9",x"000012f6",x"000012f3",
		x"000012f0",x"000012ed",x"000012e9",x"000012e6",x"000012e3",x"000012e0",x"000012dd",x"000012da",
		x"000012d7",x"000012d3",x"000012d0",x"000012cd",x"000012ca",x"000012c7",x"000012c4",x"000012c1",
		x"000012bd",x"000012ba",x"000012b7",x"000012b4",x"000012b1",x"000012ae",x"000012ab",x"000012a7",
		x"000012a4",x"000012a1",x"0000129e",x"0000129b",x"00001298",x"00001295",x"00001291",x"0000128e",
		x"0000128b",x"00001288",x"00001285",x"00001282",x"0000127f",x"0000127b",x"00001278",x"00001275",
		x"00001272",x"0000126f",x"0000126c",x"00001269",x"00001266",x"00001262",x"0000125f",x"0000125c",
		x"00001259",x"00001256",x"00001253",x"00001250",x"0000124c",x"00001249",x"00001246",x"00001243",
		x"00001240",x"0000123d",x"0000123a",x"00001237",x"00001233",x"00001230",x"0000122d",x"0000122a",
		x"00001227",x"00001224",x"00001221",x"0000121d",x"0000121a",x"00001217",x"00001214",x"00001211",
		x"0000120e",x"0000120b",x"00001207",x"00001204",x"00001201",x"000011fe",x"000011fb",x"000011f8",
		x"000011f5",x"000011f2",x"000011ee",x"000011eb",x"000011e8",x"000011e5",x"000011e2",x"000011df",
		x"000011dc",x"000011d9",x"000011d5",x"000011d2",x"000011cf",x"000011cc",x"000011c9",x"000011c6",
		x"000011c3",x"000011bf",x"000011bc",x"000011b9",x"000011b6",x"000011b3",x"000011b0",x"000011ad",
		x"000011aa",x"000011a6",x"000011a3",x"000011a0",x"0000119d",x"0000119a",x"00001197",x"00001194",
		x"00001191",x"0000118d",x"0000118a",x"00001187",x"00001184",x"00001181",x"0000117e",x"0000117b",
		x"00001178",x"00001174",x"00001171",x"0000116e",x"0000116b",x"00001168",x"00001165",x"00001162",
		x"0000115f",x"0000115b",x"00001158",x"00001155",x"00001152",x"0000114f",x"0000114c",x"00001149",
		x"00001146",x"00001142",x"0000113f",x"0000113c",x"00001139",x"00001136",x"00001133",x"00001130",
		x"0000112d",x"0000112a",x"00001126",x"00001123",x"00001120",x"0000111d",x"0000111a",x"00001117",
		x"00001114",x"00001111",x"0000110d",x"0000110a",x"00001107",x"00001104",x"00001101",x"000010fe",
		x"000010fb",x"000010f8",x"000010f5",x"000010f1",x"000010ee",x"000010eb",x"000010e8",x"000010e5",
		x"000010e2",x"000010df",x"000010dc",x"000010d9",x"000010d5",x"000010d2",x"000010cf",x"000010cc",
		x"000010c9",x"000010c6",x"000010c3",x"000010c0",x"000010bd",x"000010b9",x"000010b6",x"000010b3",
		x"000010b0",x"000010ad",x"000010aa",x"000010a7",x"000010a4",x"000010a1",x"0000109d",x"0000109a",
		x"00001097",x"00001094",x"00001091",x"0000108e",x"0000108b",x"00001088",x"00001085",x"00001082",
		x"0000107e",x"0000107b",x"00001078",x"00001075",x"00001072",x"0000106f",x"0000106c",x"00001069",
		x"00001066",x"00001062",x"0000105f",x"0000105c",x"00001059",x"00001056",x"00001053",x"00001050",
		x"0000104d",x"0000104a",x"00001047",x"00001043",x"00001040",x"0000103d",x"0000103a",x"00001037",
		x"00001034",x"00001031",x"0000102e",x"0000102b",x"00001028",x"00001025",x"00001021",x"0000101e",
		x"0000101b",x"00001018",x"00001015",x"00001012",x"0000100f",x"0000100c",x"00001009",x"00001006",
		x"00001003",x"00000fff",x"00000ffc",x"00000ff9",x"00000ff6",x"00000ff3",x"00000ff0",x"00000fed",
		x"00000fea",x"00000fe7",x"00000fe4",x"00000fe1",x"00000fdd",x"00000fda",x"00000fd7",x"00000fd4",
		x"00000fd1",x"00000fce",x"00000fcb",x"00000fc8",x"00000fc5",x"00000fc2",x"00000fbf",x"00000fbc",
		x"00000fb8",x"00000fb5",x"00000fb2",x"00000faf",x"00000fac",x"00000fa9",x"00000fa6",x"00000fa3",
		x"00000fa0",x"00000f9d",x"00000f9a",x"00000f97",x"00000f94",x"00000f90",x"00000f8d",x"00000f8a",
		x"00000f87",x"00000f84",x"00000f81",x"00000f7e",x"00000f7b",x"00000f78",x"00000f75",x"00000f72",
		x"00000f6f",x"00000f6c",x"00000f68",x"00000f65",x"00000f62",x"00000f5f",x"00000f5c",x"00000f59",
		x"00000f56",x"00000f53",x"00000f50",x"00000f4d",x"00000f4a",x"00000f47",x"00000f44",x"00000f41",
		x"00000f3e",x"00000f3a",x"00000f37",x"00000f34",x"00000f31",x"00000f2e",x"00000f2b",x"00000f28",
		x"00000f25",x"00000f22",x"00000f1f",x"00000f1c",x"00000f19",x"00000f16",x"00000f13",x"00000f10",
		x"00000f0d",x"00000f09",x"00000f06",x"00000f03",x"00000f00",x"00000efd",x"00000efa",x"00000ef7",
		x"00000ef4",x"00000ef1",x"00000eee",x"00000eeb",x"00000ee8",x"00000ee5",x"00000ee2",x"00000edf",
		x"00000edc",x"00000ed9",x"00000ed6",x"00000ed3",x"00000ecf",x"00000ecc",x"00000ec9",x"00000ec6",
		x"00000ec3",x"00000ec0",x"00000ebd",x"00000eba",x"00000eb7",x"00000eb4",x"00000eb1",x"00000eae",
		x"00000eab",x"00000ea8",x"00000ea5",x"00000ea2",x"00000e9f",x"00000e9c",x"00000e99",x"00000e96",
		x"00000e93",x"00000e90",x"00000e8d",x"00000e89",x"00000e86",x"00000e83",x"00000e80",x"00000e7d",
		x"00000e7a",x"00000e77",x"00000e74",x"00000e71",x"00000e6e",x"00000e6b",x"00000e68",x"00000e65",
		x"00000e62",x"00000e5f",x"00000e5c",x"00000e59",x"00000e56",x"00000e53",x"00000e50",x"00000e4d",
		x"00000e4a",x"00000e47",x"00000e44",x"00000e41",x"00000e3e",x"00000e3b",x"00000e38",x"00000e35",
		x"00000e32",x"00000e2f",x"00000e2c",x"00000e29",x"00000e26",x"00000e22",x"00000e1f",x"00000e1c",
		x"00000e19",x"00000e16",x"00000e13",x"00000e10",x"00000e0d",x"00000e0a",x"00000e07",x"00000e04",
		x"00000e01",x"00000dfe",x"00000dfb",x"00000df8",x"00000df5",x"00000df2",x"00000def",x"00000dec",
		x"00000de9",x"00000de6",x"00000de3",x"00000de0",x"00000ddd",x"00000dda",x"00000dd7",x"00000dd4",
		x"00000dd1",x"00000dce",x"00000dcb",x"00000dc8",x"00000dc5",x"00000dc2",x"00000dbf",x"00000dbc",
		x"00000db9",x"00000db6",x"00000db3",x"00000db0",x"00000dad",x"00000daa",x"00000da7",x"00000da4",
		x"00000da1",x"00000d9e",x"00000d9b",x"00000d98",x"00000d95",x"00000d92",x"00000d8f",x"00000d8c",
		x"00000d89",x"00000d86",x"00000d83",x"00000d80",x"00000d7d",x"00000d7a",x"00000d77",x"00000d74",
		x"00000d71",x"00000d6e",x"00000d6b",x"00000d68",x"00000d65",x"00000d62",x"00000d5f",x"00000d5c",
		x"00000d59",x"00000d56",x"00000d54",x"00000d51",x"00000d4e",x"00000d4b",x"00000d48",x"00000d45",
		x"00000d42",x"00000d3f",x"00000d3c",x"00000d39",x"00000d36",x"00000d33",x"00000d30",x"00000d2d",
		x"00000d2a",x"00000d27",x"00000d24",x"00000d21",x"00000d1e",x"00000d1b",x"00000d18",x"00000d15",
		x"00000d12",x"00000d0f",x"00000d0c",x"00000d09",x"00000d06",x"00000d03",x"00000d00",x"00000cfd",
		x"00000cfa",x"00000cf7",x"00000cf4",x"00000cf2",x"00000cef",x"00000cec",x"00000ce9",x"00000ce6",
		x"00000ce3",x"00000ce0",x"00000cdd",x"00000cda",x"00000cd7",x"00000cd4",x"00000cd1",x"00000cce",
		x"00000ccb",x"00000cc8",x"00000cc5",x"00000cc2",x"00000cbf",x"00000cbc",x"00000cb9",x"00000cb7",
		x"00000cb4",x"00000cb1",x"00000cae",x"00000cab",x"00000ca8",x"00000ca5",x"00000ca2",x"00000c9f",
		x"00000c9c",x"00000c99",x"00000c96",x"00000c93",x"00000c90",x"00000c8d",x"00000c8a",x"00000c88",
		x"00000c85",x"00000c82",x"00000c7f",x"00000c7c",x"00000c79",x"00000c76",x"00000c73",x"00000c70",
		x"00000c6d",x"00000c6a",x"00000c67",x"00000c64",x"00000c61",x"00000c5f",x"00000c5c",x"00000c59",
		x"00000c56",x"00000c53",x"00000c50",x"00000c4d",x"00000c4a",x"00000c47",x"00000c44",x"00000c41",
		x"00000c3e",x"00000c3b",x"00000c39",x"00000c36",x"00000c33",x"00000c30",x"00000c2d",x"00000c2a",
		x"00000c27",x"00000c24",x"00000c21",x"00000c1e",x"00000c1b",x"00000c19",x"00000c16",x"00000c13",
		x"00000c10",x"00000c0d",x"00000c0a",x"00000c07",x"00000c04",x"00000c01",x"00000bfe",x"00000bfc",
		x"00000bf9",x"00000bf6",x"00000bf3",x"00000bf0",x"00000bed",x"00000bea",x"00000be7",x"00000be4",
		x"00000be2",x"00000bdf",x"00000bdc",x"00000bd9",x"00000bd6",x"00000bd3",x"00000bd0",x"00000bcd",
		x"00000bca",x"00000bc8",x"00000bc5",x"00000bc2",x"00000bbf",x"00000bbc",x"00000bb9",x"00000bb6",
		x"00000bb3",x"00000bb0",x"00000bae",x"00000bab",x"00000ba8",x"00000ba5",x"00000ba2",x"00000b9f",
		x"00000b9c",x"00000b99",x"00000b97",x"00000b94",x"00000b91",x"00000b8e",x"00000b8b",x"00000b88",
		x"00000b85",x"00000b83",x"00000b80",x"00000b7d",x"00000b7a",x"00000b77",x"00000b74",x"00000b71",
		x"00000b6e",x"00000b6c",x"00000b69",x"00000b66",x"00000b63",x"00000b60",x"00000b5d",x"00000b5b",
		x"00000b58",x"00000b55",x"00000b52",x"00000b4f",x"00000b4c",x"00000b49",x"00000b47",x"00000b44",
		x"00000b41",x"00000b3e",x"00000b3b",x"00000b38",x"00000b35",x"00000b33",x"00000b30",x"00000b2d",
		x"00000b2a",x"00000b27",x"00000b24",x"00000b22",x"00000b1f",x"00000b1c",x"00000b19",x"00000b16",
		x"00000b13",x"00000b11",x"00000b0e",x"00000b0b",x"00000b08",x"00000b05",x"00000b02",x"00000b00",
		x"00000afd",x"00000afa",x"00000af7",x"00000af4",x"00000af2",x"00000aef",x"00000aec",x"00000ae9",
		x"00000ae6",x"00000ae3",x"00000ae1",x"00000ade",x"00000adb",x"00000ad8",x"00000ad5",x"00000ad3",
		x"00000ad0",x"00000acd",x"00000aca",x"00000ac7",x"00000ac4",x"00000ac2",x"00000abf",x"00000abc",
		x"00000ab9",x"00000ab6",x"00000ab4",x"00000ab1",x"00000aae",x"00000aab",x"00000aa8",x"00000aa6",
		x"00000aa3",x"00000aa0",x"00000a9d",x"00000a9a",x"00000a98",x"00000a95",x"00000a92",x"00000a8f",
		x"00000a8c",x"00000a8a",x"00000a87",x"00000a84",x"00000a81",x"00000a7f",x"00000a7c",x"00000a79",
		x"00000a76",x"00000a73",x"00000a71",x"00000a6e",x"00000a6b",x"00000a68",x"00000a66",x"00000a63",
		x"00000a60",x"00000a5d",x"00000a5a",x"00000a58",x"00000a55",x"00000a52",x"00000a4f",x"00000a4d",
		x"00000a4a",x"00000a47",x"00000a44",x"00000a42",x"00000a3f",x"00000a3c",x"00000a39",x"00000a36",
		x"00000a34",x"00000a31",x"00000a2e",x"00000a2b",x"00000a29",x"00000a26",x"00000a23",x"00000a20",
		x"00000a1e",x"00000a1b",x"00000a18",x"00000a15",x"00000a13",x"00000a10",x"00000a0d",x"00000a0a",
		x"00000a08",x"00000a05",x"00000a02",x"000009ff",x"000009fd",x"000009fa",x"000009f7",x"000009f4",
		x"000009f2",x"000009ef",x"000009ec",x"000009ea",x"000009e7",x"000009e4",x"000009e1",x"000009df",
		x"000009dc",x"000009d9",x"000009d6",x"000009d4",x"000009d1",x"000009ce",x"000009cb",x"000009c9",
		x"000009c6",x"000009c3",x"000009c1",x"000009be",x"000009bb",x"000009b8",x"000009b6",x"000009b3",
		x"000009b0",x"000009ae",x"000009ab",x"000009a8",x"000009a5",x"000009a3",x"000009a0",x"0000099d",
		x"0000099b",x"00000998",x"00000995",x"00000993",x"00000990",x"0000098d",x"0000098a",x"00000988",
		x"00000985",x"00000982",x"00000980",x"0000097d",x"0000097a",x"00000978",x"00000975",x"00000972",
		x"0000096f",x"0000096d",x"0000096a",x"00000967",x"00000965",x"00000962",x"0000095f",x"0000095d",
		x"0000095a",x"00000957",x"00000955",x"00000952",x"0000094f",x"0000094d",x"0000094a",x"00000947",
		x"00000945",x"00000942",x"0000093f",x"0000093d",x"0000093a",x"00000937",x"00000935",x"00000932",
		x"0000092f",x"0000092d",x"0000092a",x"00000927",x"00000925",x"00000922",x"0000091f",x"0000091d",
		x"0000091a",x"00000917",x"00000915",x"00000912",x"0000090f",x"0000090d",x"0000090a",x"00000907",
		x"00000905",x"00000902",x"000008ff",x"000008fd",x"000008fa",x"000008f7",x"000008f5",x"000008f2",
		x"000008f0",x"000008ed",x"000008ea",x"000008e8",x"000008e5",x"000008e2",x"000008e0",x"000008dd",
		x"000008da",x"000008d8",x"000008d5",x"000008d3",x"000008d0",x"000008cd",x"000008cb",x"000008c8",
		x"000008c5",x"000008c3",x"000008c0",x"000008be",x"000008bb",x"000008b8",x"000008b6",x"000008b3",
		x"000008b1",x"000008ae",x"000008ab",x"000008a9",x"000008a6",x"000008a3",x"000008a1",x"0000089e",
		x"0000089c",x"00000899",x"00000896",x"00000894",x"00000891",x"0000088f",x"0000088c",x"00000889",
		x"00000887",x"00000884",x"00000882",x"0000087f",x"0000087c",x"0000087a",x"00000877",x"00000875",
		x"00000872",x"00000870",x"0000086d",x"0000086a",x"00000868",x"00000865",x"00000863",x"00000860",
		x"0000085d",x"0000085b",x"00000858",x"00000856",x"00000853",x"00000851",x"0000084e",x"0000084b",
		x"00000849",x"00000846",x"00000844",x"00000841",x"0000083f",x"0000083c",x"00000839",x"00000837",
		x"00000834",x"00000832",x"0000082f",x"0000082d",x"0000082a",x"00000828",x"00000825",x"00000822",
		x"00000820",x"0000081d",x"0000081b",x"00000818",x"00000816",x"00000813",x"00000811",x"0000080e",
		x"0000080c",x"00000809",x"00000806",x"00000804",x"00000801",x"000007ff",x"000007fc",x"000007fa",
		x"000007f7",x"000007f5",x"000007f2",x"000007f0",x"000007ed",x"000007eb",x"000007e8",x"000007e6",
		x"000007e3",x"000007e1",x"000007de",x"000007db",x"000007d9",x"000007d6",x"000007d4",x"000007d1",
		x"000007cf",x"000007cc",x"000007ca",x"000007c7",x"000007c5",x"000007c2",x"000007c0",x"000007bd",
		x"000007bb",x"000007b8",x"000007b6",x"000007b3",x"000007b1",x"000007ae",x"000007ac",x"000007a9",
		x"000007a7",x"000007a4",x"000007a2",x"0000079f",x"0000079d",x"0000079a",x"00000798",x"00000795",
		x"00000793",x"00000790",x"0000078e",x"0000078b",x"00000789",x"00000787",x"00000784",x"00000782",
		x"0000077f",x"0000077d",x"0000077a",x"00000778",x"00000775",x"00000773",x"00000770",x"0000076e",
		x"0000076b",x"00000769",x"00000766",x"00000764",x"00000761",x"0000075f",x"0000075d",x"0000075a",
		x"00000758",x"00000755",x"00000753",x"00000750",x"0000074e",x"0000074b",x"00000749",x"00000747",
		x"00000744",x"00000742",x"0000073f",x"0000073d",x"0000073a",x"00000738",x"00000735",x"00000733",
		x"00000731",x"0000072e",x"0000072c",x"00000729",x"00000727",x"00000724",x"00000722",x"00000720",
		x"0000071d",x"0000071b",x"00000718",x"00000716",x"00000713",x"00000711",x"0000070f",x"0000070c",
		x"0000070a",x"00000707",x"00000705",x"00000702",x"00000700",x"000006fe",x"000006fb",x"000006f9",
		x"000006f6",x"000006f4",x"000006f2",x"000006ef",x"000006ed",x"000006ea",x"000006e8",x"000006e6",
		x"000006e3",x"000006e1",x"000006de",x"000006dc",x"000006da",x"000006d7",x"000006d5",x"000006d3",
		x"000006d0",x"000006ce",x"000006cb",x"000006c9",x"000006c7",x"000006c4",x"000006c2",x"000006bf",
		x"000006bd",x"000006bb",x"000006b8",x"000006b6",x"000006b4",x"000006b1",x"000006af",x"000006ad",
		x"000006aa",x"000006a8",x"000006a5",x"000006a3",x"000006a1",x"0000069e",x"0000069c",x"0000069a",
		x"00000697",x"00000695",x"00000693",x"00000690",x"0000068e",x"0000068c",x"00000689",x"00000687",
		x"00000684",x"00000682",x"00000680",x"0000067d",x"0000067b",x"00000679",x"00000676",x"00000674",
		x"00000672",x"0000066f",x"0000066d",x"0000066b",x"00000668",x"00000666",x"00000664",x"00000662",
		x"0000065f",x"0000065d",x"0000065b",x"00000658",x"00000656",x"00000654",x"00000651",x"0000064f",
		x"0000064d",x"0000064a",x"00000648",x"00000646",x"00000643",x"00000641",x"0000063f",x"0000063d",
		x"0000063a",x"00000638",x"00000636",x"00000633",x"00000631",x"0000062f",x"0000062c",x"0000062a",
		x"00000628",x"00000626",x"00000623",x"00000621",x"0000061f",x"0000061c",x"0000061a",x"00000618",
		x"00000616",x"00000613",x"00000611",x"0000060f",x"0000060c",x"0000060a",x"00000608",x"00000606",
		x"00000603",x"00000601",x"000005ff",x"000005fd",x"000005fa",x"000005f8",x"000005f6",x"000005f4",
		x"000005f1",x"000005ef",x"000005ed",x"000005eb",x"000005e8",x"000005e6",x"000005e4",x"000005e2",
		x"000005df",x"000005dd",x"000005db",x"000005d9",x"000005d6",x"000005d4",x"000005d2",x"000005d0",
		x"000005cd",x"000005cb",x"000005c9",x"000005c7",x"000005c4",x"000005c2",x"000005c0",x"000005be",
		x"000005bc",x"000005b9",x"000005b7",x"000005b5",x"000005b3",x"000005b0",x"000005ae",x"000005ac",
		x"000005aa",x"000005a8",x"000005a5",x"000005a3",x"000005a1",x"0000059f",x"0000059d",x"0000059a",
		x"00000598",x"00000596",x"00000594",x"00000592",x"0000058f",x"0000058d",x"0000058b",x"00000589",
		x"00000587",x"00000584",x"00000582",x"00000580",x"0000057e",x"0000057c",x"00000579",x"00000577",
		x"00000575",x"00000573",x"00000571",x"0000056f",x"0000056c",x"0000056a",x"00000568",x"00000566",
		x"00000564",x"00000562",x"0000055f",x"0000055d",x"0000055b",x"00000559",x"00000557",x"00000555",
		x"00000552",x"00000550",x"0000054e",x"0000054c",x"0000054a",x"00000548",x"00000546",x"00000543",
		x"00000541",x"0000053f",x"0000053d",x"0000053b",x"00000539",x"00000537",x"00000534",x"00000532",
		x"00000530",x"0000052e",x"0000052c",x"0000052a",x"00000528",x"00000525",x"00000523",x"00000521",
		x"0000051f",x"0000051d",x"0000051b",x"00000519",x"00000517",x"00000515",x"00000512",x"00000510",
		x"0000050e",x"0000050c",x"0000050a",x"00000508",x"00000506",x"00000504",x"00000502",x"000004ff",
		x"000004fd",x"000004fb",x"000004f9",x"000004f7",x"000004f5",x"000004f3",x"000004f1",x"000004ef",
		x"000004ed",x"000004eb",x"000004e8",x"000004e6",x"000004e4",x"000004e2",x"000004e0",x"000004de",
		x"000004dc",x"000004da",x"000004d8",x"000004d6",x"000004d4",x"000004d2",x"000004d0",x"000004cd",
		x"000004cb",x"000004c9",x"000004c7",x"000004c5",x"000004c3",x"000004c1",x"000004bf",x"000004bd",
		x"000004bb",x"000004b9",x"000004b7",x"000004b5",x"000004b3",x"000004b1",x"000004af",x"000004ad",
		x"000004ab",x"000004a9",x"000004a7",x"000004a5",x"000004a2",x"000004a0",x"0000049e",x"0000049c",
		x"0000049a",x"00000498",x"00000496",x"00000494",x"00000492",x"00000490",x"0000048e",x"0000048c",
		x"0000048a",x"00000488",x"00000486",x"00000484",x"00000482",x"00000480",x"0000047e",x"0000047c",
		x"0000047a",x"00000478",x"00000476",x"00000474",x"00000472",x"00000470",x"0000046e",x"0000046c",
		x"0000046a",x"00000468",x"00000466",x"00000464",x"00000462",x"00000460",x"0000045e",x"0000045c",
		x"0000045a",x"00000458",x"00000456",x"00000454",x"00000452",x"00000450",x"0000044e",x"0000044d",
		x"0000044b",x"00000449",x"00000447",x"00000445",x"00000443",x"00000441",x"0000043f",x"0000043d",
		x"0000043b",x"00000439",x"00000437",x"00000435",x"00000433",x"00000431",x"0000042f",x"0000042d",
		x"0000042b",x"00000429",x"00000427",x"00000425",x"00000424",x"00000422",x"00000420",x"0000041e",
		x"0000041c",x"0000041a",x"00000418",x"00000416",x"00000414",x"00000412",x"00000410",x"0000040e",
		x"0000040c",x"0000040b",x"00000409",x"00000407",x"00000405",x"00000403",x"00000401",x"000003ff",
		x"000003fd",x"000003fb",x"000003f9",x"000003f7",x"000003f6",x"000003f4",x"000003f2",x"000003f0",
		x"000003ee",x"000003ec",x"000003ea",x"000003e8",x"000003e6",x"000003e5",x"000003e3",x"000003e1",
		x"000003df",x"000003dd",x"000003db",x"000003d9",x"000003d7",x"000003d6",x"000003d4",x"000003d2",
		x"000003d0",x"000003ce",x"000003cc",x"000003ca",x"000003c9",x"000003c7",x"000003c5",x"000003c3",
		x"000003c1",x"000003bf",x"000003bd",x"000003bc",x"000003ba",x"000003b8",x"000003b6",x"000003b4",
		x"000003b2",x"000003b1",x"000003af",x"000003ad",x"000003ab",x"000003a9",x"000003a7",x"000003a6",
		x"000003a4",x"000003a2",x"000003a0",x"0000039e",x"0000039c",x"0000039b",x"00000399",x"00000397",
		x"00000395",x"00000393",x"00000391",x"00000390",x"0000038e",x"0000038c",x"0000038a",x"00000388",
		x"00000387",x"00000385",x"00000383",x"00000381",x"0000037f",x"0000037e",x"0000037c",x"0000037a",
		x"00000378",x"00000377",x"00000375",x"00000373",x"00000371",x"0000036f",x"0000036e",x"0000036c",
		x"0000036a",x"00000368",x"00000367",x"00000365",x"00000363",x"00000361",x"0000035f",x"0000035e",
		x"0000035c",x"0000035a",x"00000358",x"00000357",x"00000355",x"00000353",x"00000351",x"00000350",
		x"0000034e",x"0000034c",x"0000034a",x"00000349",x"00000347",x"00000345",x"00000343",x"00000342",
		x"00000340",x"0000033e",x"0000033c",x"0000033b",x"00000339",x"00000337",x"00000336",x"00000334",
		x"00000332",x"00000330",x"0000032f",x"0000032d",x"0000032b",x"0000032a",x"00000328",x"00000326",
		x"00000324",x"00000323",x"00000321",x"0000031f",x"0000031e",x"0000031c",x"0000031a",x"00000318",
		x"00000317",x"00000315",x"00000313",x"00000312",x"00000310",x"0000030e",x"0000030d",x"0000030b",
		x"00000309",x"00000308",x"00000306",x"00000304",x"00000303",x"00000301",x"000002ff",x"000002fe",
		x"000002fc",x"000002fa",x"000002f9",x"000002f7",x"000002f5",x"000002f4",x"000002f2",x"000002f0",
		x"000002ef",x"000002ed",x"000002eb",x"000002ea",x"000002e8",x"000002e6",x"000002e5",x"000002e3",
		x"000002e1",x"000002e0",x"000002de",x"000002dc",x"000002db",x"000002d9",x"000002d8",x"000002d6",
		x"000002d4",x"000002d3",x"000002d1",x"000002cf",x"000002ce",x"000002cc",x"000002cb",x"000002c9",
		x"000002c7",x"000002c6",x"000002c4",x"000002c2",x"000002c1",x"000002bf",x"000002be",x"000002bc",
		x"000002ba",x"000002b9",x"000002b7",x"000002b6",x"000002b4",x"000002b2",x"000002b1",x"000002af",
		x"000002ae",x"000002ac",x"000002aa",x"000002a9",x"000002a7",x"000002a6",x"000002a4",x"000002a3",
		x"000002a1",x"0000029f",x"0000029e",x"0000029c",x"0000029b",x"00000299",x"00000298",x"00000296",
		x"00000294",x"00000293",x"00000291",x"00000290",x"0000028e",x"0000028d",x"0000028b",x"0000028a",
		x"00000288",x"00000287",x"00000285",x"00000283",x"00000282",x"00000280",x"0000027f",x"0000027d",
		x"0000027c",x"0000027a",x"00000279",x"00000277",x"00000276",x"00000274",x"00000273",x"00000271",
		x"00000270",x"0000026e",x"0000026c",x"0000026b",x"00000269",x"00000268",x"00000266",x"00000265",
		x"00000263",x"00000262",x"00000260",x"0000025f",x"0000025d",x"0000025c",x"0000025a",x"00000259",
		x"00000257",x"00000256",x"00000254",x"00000253",x"00000251",x"00000250",x"0000024f",x"0000024d",
		x"0000024c",x"0000024a",x"00000249",x"00000247",x"00000246",x"00000244",x"00000243",x"00000241",
		x"00000240",x"0000023e",x"0000023d",x"0000023b",x"0000023a",x"00000238",x"00000237",x"00000236",
		x"00000234",x"00000233",x"00000231",x"00000230",x"0000022e",x"0000022d",x"0000022b",x"0000022a",
		x"00000229",x"00000227",x"00000226",x"00000224",x"00000223",x"00000221",x"00000220",x"0000021f",
		x"0000021d",x"0000021c",x"0000021a",x"00000219",x"00000217",x"00000216",x"00000215",x"00000213",
		x"00000212",x"00000210",x"0000020f",x"0000020e",x"0000020c",x"0000020b",x"00000209",x"00000208",
		x"00000207",x"00000205",x"00000204",x"00000202",x"00000201",x"00000200",x"000001fe",x"000001fd",
		x"000001fc",x"000001fa",x"000001f9",x"000001f7",x"000001f6",x"000001f5",x"000001f3",x"000001f2",
		x"000001f1",x"000001ef",x"000001ee",x"000001ec",x"000001eb",x"000001ea",x"000001e8",x"000001e7",
		x"000001e6",x"000001e4",x"000001e3",x"000001e2",x"000001e0",x"000001df",x"000001de",x"000001dc",
		x"000001db",x"000001da",x"000001d8",x"000001d7",x"000001d6",x"000001d4",x"000001d3",x"000001d2",
		x"000001d0",x"000001cf",x"000001ce",x"000001cc",x"000001cb",x"000001ca",x"000001c8",x"000001c7",
		x"000001c6",x"000001c4",x"000001c3",x"000001c2",x"000001c1",x"000001bf",x"000001be",x"000001bd",
		x"000001bb",x"000001ba",x"000001b9",x"000001b8",x"000001b6",x"000001b5",x"000001b4",x"000001b2",
		x"000001b1",x"000001b0",x"000001af",x"000001ad",x"000001ac",x"000001ab",x"000001a9",x"000001a8",
		x"000001a7",x"000001a6",x"000001a4",x"000001a3",x"000001a2",x"000001a1",x"0000019f",x"0000019e",
		x"0000019d",x"0000019c",x"0000019a",x"00000199",x"00000198",x"00000197",x"00000195",x"00000194",
		x"00000193",x"00000192",x"00000190",x"0000018f",x"0000018e",x"0000018d",x"0000018c",x"0000018a",
		x"00000189",x"00000188",x"00000187",x"00000185",x"00000184",x"00000183",x"00000182",x"00000181",
		x"0000017f",x"0000017e",x"0000017d",x"0000017c",x"0000017b",x"00000179",x"00000178",x"00000177",
		x"00000176",x"00000175",x"00000173",x"00000172",x"00000171",x"00000170",x"0000016f",x"0000016d",
		x"0000016c",x"0000016b",x"0000016a",x"00000169",x"00000168",x"00000166",x"00000165",x"00000164",
		x"00000163",x"00000162",x"00000161",x"0000015f",x"0000015e",x"0000015d",x"0000015c",x"0000015b",
		x"0000015a",x"00000159",x"00000157",x"00000156",x"00000155",x"00000154",x"00000153",x"00000152",
		x"00000151",x"0000014f",x"0000014e",x"0000014d",x"0000014c",x"0000014b",x"0000014a",x"00000149",
		x"00000148",x"00000146",x"00000145",x"00000144",x"00000143",x"00000142",x"00000141",x"00000140",
		x"0000013f",x"0000013e",x"0000013c",x"0000013b",x"0000013a",x"00000139",x"00000138",x"00000137",
		x"00000136",x"00000135",x"00000134",x"00000133",x"00000132",x"00000130",x"0000012f",x"0000012e",
		x"0000012d",x"0000012c",x"0000012b",x"0000012a",x"00000129",x"00000128",x"00000127",x"00000126",
		x"00000125",x"00000124",x"00000123",x"00000122",x"00000121",x"0000011f",x"0000011e",x"0000011d",
		x"0000011c",x"0000011b",x"0000011a",x"00000119",x"00000118",x"00000117",x"00000116",x"00000115",
		x"00000114",x"00000113",x"00000112",x"00000111",x"00000110",x"0000010f",x"0000010e",x"0000010d",
		x"0000010c",x"0000010b",x"0000010a",x"00000109",x"00000108",x"00000107",x"00000106",x"00000105",
		x"00000104",x"00000103",x"00000102",x"00000101",x"00000100",x"000000ff",x"000000fe",x"000000fd",
		x"000000fc",x"000000fb",x"000000fa",x"000000f9",x"000000f8",x"000000f7",x"000000f6",x"000000f5",
		x"000000f4",x"000000f3",x"000000f2",x"000000f1",x"000000f0",x"000000ef",x"000000ee",x"000000ed",
		x"000000ec",x"000000eb",x"000000ea",x"000000e9",x"000000e9",x"000000e8",x"000000e7",x"000000e6",
		x"000000e5",x"000000e4",x"000000e3",x"000000e2",x"000000e1",x"000000e0",x"000000df",x"000000de",
		x"000000dd",x"000000dc",x"000000db",x"000000db",x"000000da",x"000000d9",x"000000d8",x"000000d7",
		x"000000d6",x"000000d5",x"000000d4",x"000000d3",x"000000d2",x"000000d1",x"000000d1",x"000000d0",
		x"000000cf",x"000000ce",x"000000cd",x"000000cc",x"000000cb",x"000000ca",x"000000c9",x"000000c9",
		x"000000c8",x"000000c7",x"000000c6",x"000000c5",x"000000c4",x"000000c3",x"000000c2",x"000000c2",
		x"000000c1",x"000000c0",x"000000bf",x"000000be",x"000000bd",x"000000bc",x"000000bc",x"000000bb",
		x"000000ba",x"000000b9",x"000000b8",x"000000b7",x"000000b6",x"000000b6",x"000000b5",x"000000b4",
		x"000000b3",x"000000b2",x"000000b1",x"000000b1",x"000000b0",x"000000af",x"000000ae",x"000000ad",
		x"000000ad",x"000000ac",x"000000ab",x"000000aa",x"000000a9",x"000000a8",x"000000a8",x"000000a7",
		x"000000a6",x"000000a5",x"000000a4",x"000000a4",x"000000a3",x"000000a2",x"000000a1",x"000000a0",
		x"000000a0",x"0000009f",x"0000009e",x"0000009d",x"0000009d",x"0000009c",x"0000009b",x"0000009a",
		x"00000099",x"00000099",x"00000098",x"00000097",x"00000096",x"00000096",x"00000095",x"00000094",
		x"00000093",x"00000093",x"00000092",x"00000091",x"00000090",x"00000090",x"0000008f",x"0000008e",
		x"0000008d",x"0000008d",x"0000008c",x"0000008b",x"0000008a",x"0000008a",x"00000089",x"00000088",
		x"00000087",x"00000087",x"00000086",x"00000085",x"00000085",x"00000084",x"00000083",x"00000082",
		x"00000082",x"00000081",x"00000080",x"00000080",x"0000007f",x"0000007e",x"0000007d",x"0000007d",
		x"0000007c",x"0000007b",x"0000007b",x"0000007a",x"00000079",x"00000079",x"00000078",x"00000077",
		x"00000077",x"00000076",x"00000075",x"00000075",x"00000074",x"00000073",x"00000073",x"00000072",
		x"00000071",x"00000071",x"00000070",x"0000006f",x"0000006f",x"0000006e",x"0000006d",x"0000006d",
		x"0000006c",x"0000006b",x"0000006b",x"0000006a",x"00000069",x"00000069",x"00000068",x"00000067",
		x"00000067",x"00000066",x"00000066",x"00000065",x"00000064",x"00000064",x"00000063",x"00000062",
		x"00000062",x"00000061",x"00000061",x"00000060",x"0000005f",x"0000005f",x"0000005e",x"0000005e",
		x"0000005d",x"0000005c",x"0000005c",x"0000005b",x"0000005b",x"0000005a",x"00000059",x"00000059",
		x"00000058",x"00000058",x"00000057",x"00000056",x"00000056",x"00000055",x"00000055",x"00000054",
		x"00000054",x"00000053",x"00000052",x"00000052",x"00000051",x"00000051",x"00000050",x"00000050",
		x"0000004f",x"0000004e",x"0000004e",x"0000004d",x"0000004d",x"0000004c",x"0000004c",x"0000004b",
		x"0000004b",x"0000004a",x"0000004a",x"00000049",x"00000048",x"00000048",x"00000047",x"00000047",
		x"00000046",x"00000046",x"00000045",x"00000045",x"00000044",x"00000044",x"00000043",x"00000043",
		x"00000042",x"00000042",x"00000041",x"00000041",x"00000040",x"00000040",x"0000003f",x"0000003f",
		x"0000003e",x"0000003e",x"0000003d",x"0000003d",x"0000003c",x"0000003c",x"0000003b",x"0000003b",
		x"0000003a",x"0000003a",x"00000039",x"00000039",x"00000038",x"00000038",x"00000037",x"00000037",
		x"00000037",x"00000036",x"00000036",x"00000035",x"00000035",x"00000034",x"00000034",x"00000033",
		x"00000033",x"00000032",x"00000032",x"00000032",x"00000031",x"00000031",x"00000030",x"00000030",
		x"0000002f",x"0000002f",x"0000002f",x"0000002e",x"0000002e",x"0000002d",x"0000002d",x"0000002c",
		x"0000002c",x"0000002c",x"0000002b",x"0000002b",x"0000002a",x"0000002a",x"0000002a",x"00000029",
		x"00000029",x"00000028",x"00000028",x"00000028",x"00000027",x"00000027",x"00000026",x"00000026",
		x"00000026",x"00000025",x"00000025",x"00000024",x"00000024",x"00000024",x"00000023",x"00000023",
		x"00000023",x"00000022",x"00000022",x"00000021",x"00000021",x"00000021",x"00000020",x"00000020",
		x"00000020",x"0000001f",x"0000001f",x"0000001f",x"0000001e",x"0000001e",x"0000001e",x"0000001d",
		x"0000001d",x"0000001d",x"0000001c",x"0000001c",x"0000001c",x"0000001b",x"0000001b",x"0000001b",
		x"0000001a",x"0000001a",x"0000001a",x"00000019",x"00000019",x"00000019",x"00000018",x"00000018",
		x"00000018",x"00000017",x"00000017",x"00000017",x"00000017",x"00000016",x"00000016",x"00000016",
		x"00000015",x"00000015",x"00000015",x"00000015",x"00000014",x"00000014",x"00000014",x"00000013",
		x"00000013",x"00000013",x"00000013",x"00000012",x"00000012",x"00000012",x"00000012",x"00000011",
		x"00000011",x"00000011",x"00000010",x"00000010",x"00000010",x"00000010",x"0000000f",x"0000000f",
		x"0000000f",x"0000000f",x"0000000f",x"0000000e",x"0000000e",x"0000000e",x"0000000e",x"0000000d",
		x"0000000d",x"0000000d",x"0000000d",x"0000000c",x"0000000c",x"0000000c",x"0000000c",x"0000000c",
		x"0000000b",x"0000000b",x"0000000b",x"0000000b",x"0000000b",x"0000000a",x"0000000a",x"0000000a",
		x"0000000a",x"0000000a",x"00000009",x"00000009",x"00000009",x"00000009",x"00000009",x"00000008",
		x"00000008",x"00000008",x"00000008",x"00000008",x"00000008",x"00000007",x"00000007",x"00000007",
		x"00000007",x"00000007",x"00000007",x"00000006",x"00000006",x"00000006",x"00000006",x"00000006",
		x"00000006",x"00000005",x"00000005",x"00000005",x"00000005",x"00000005",x"00000005",x"00000005",
		x"00000004",x"00000004",x"00000004",x"00000004",x"00000004",x"00000004",x"00000004",x"00000004",
		x"00000003",x"00000003",x"00000003",x"00000003",x"00000003",x"00000003",x"00000003",x"00000003",
		x"00000003",x"00000002",x"00000002",x"00000002",x"00000002",x"00000002",x"00000002",x"00000002",
		x"00000002",x"00000002",x"00000002",x"00000002",x"00000002",x"00000001",x"00000001",x"00000001",
		x"00000001",x"00000001",x"00000001",x"00000001",x"00000001",x"00000001",x"00000001",x"00000001",
		x"00000001",x"00000001",x"00000001",x"00000001",x"00000001",x"00000000",x"00000000",x"00000000",
		x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",
		x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",
		x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",
		x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",
		x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",x"00000000",
		x"00000000",x"00000000",x"00000001",x"00000001",x"00000001",x"00000001",x"00000001",x"00000001",
		x"00000001",x"00000001",x"00000001",x"00000001",x"00000001",x"00000001",x"00000001",x"00000001",
		x"00000001",x"00000001",x"00000001",x"00000002",x"00000002",x"00000002",x"00000002",x"00000002",
		x"00000002",x"00000002",x"00000002",x"00000002",x"00000002",x"00000002",x"00000003",x"00000003",
		x"00000003",x"00000003",x"00000003",x"00000003",x"00000003",x"00000003",x"00000003",x"00000004",
		x"00000004",x"00000004",x"00000004",x"00000004",x"00000004",x"00000004",x"00000004",x"00000005",
		x"00000005",x"00000005",x"00000005",x"00000005",x"00000005",x"00000005",x"00000006",x"00000006",
		x"00000006",x"00000006",x"00000006",x"00000006",x"00000006",x"00000007",x"00000007",x"00000007",
		x"00000007",x"00000007",x"00000007",x"00000008",x"00000008",x"00000008",x"00000008",x"00000008",
		x"00000008",x"00000009",x"00000009",x"00000009",x"00000009",x"00000009",x"0000000a",x"0000000a",
		x"0000000a",x"0000000a",x"0000000a",x"0000000b",x"0000000b",x"0000000b",x"0000000b",x"0000000b",
		x"0000000c",x"0000000c",x"0000000c",x"0000000c",x"0000000d",x"0000000d",x"0000000d",x"0000000d",
		x"0000000d",x"0000000e",x"0000000e",x"0000000e",x"0000000e",x"0000000f",x"0000000f",x"0000000f",
		x"0000000f",x"00000010",x"00000010",x"00000010",x"00000010",x"00000011",x"00000011",x"00000011",
		x"00000011",x"00000012",x"00000012",x"00000012",x"00000012",x"00000013",x"00000013",x"00000013",
		x"00000014",x"00000014",x"00000014",x"00000014",x"00000015",x"00000015",x"00000015",x"00000016",
		x"00000016",x"00000016",x"00000016",x"00000017",x"00000017",x"00000017",x"00000018",x"00000018",
		x"00000018",x"00000019",x"00000019",x"00000019",x"00000019",x"0000001a",x"0000001a",x"0000001a",
		x"0000001b",x"0000001b",x"0000001b",x"0000001c",x"0000001c",x"0000001c",x"0000001d",x"0000001d",
		x"0000001d",x"0000001e",x"0000001e",x"0000001e",x"0000001f",x"0000001f",x"00000020",x"00000020",
		x"00000020",x"00000021",x"00000021",x"00000021",x"00000022",x"00000022",x"00000022",x"00000023",
		x"00000023",x"00000024",x"00000024",x"00000024",x"00000025",x"00000025",x"00000025",x"00000026",
		x"00000026",x"00000027",x"00000027",x"00000027",x"00000028",x"00000028",x"00000029",x"00000029",
		x"00000029",x"0000002a",x"0000002a",x"0000002b",x"0000002b",x"0000002b",x"0000002c",x"0000002c",
		x"0000002d",x"0000002d",x"0000002d",x"0000002e",x"0000002e",x"0000002f",x"0000002f",x"00000030",
		x"00000030",x"00000030",x"00000031",x"00000031",x"00000032",x"00000032",x"00000033",x"00000033",
		x"00000034",x"00000034",x"00000034",x"00000035",x"00000035",x"00000036",x"00000036",x"00000037",
		x"00000037",x"00000038",x"00000038",x"00000039",x"00000039",x"0000003a",x"0000003a",x"0000003b",
		x"0000003b",x"0000003b",x"0000003c",x"0000003c",x"0000003d",x"0000003d",x"0000003e",x"0000003e",
		x"0000003f",x"0000003f",x"00000040",x"00000040",x"00000041",x"00000041",x"00000042",x"00000042",
		x"00000043",x"00000043",x"00000044",x"00000045",x"00000045",x"00000046",x"00000046",x"00000047",
		x"00000047",x"00000048",x"00000048",x"00000049",x"00000049",x"0000004a",x"0000004a",x"0000004b",
		x"0000004b",x"0000004c",x"0000004d",x"0000004d",x"0000004e",x"0000004e",x"0000004f",x"0000004f",
		x"00000050",x"00000050",x"00000051",x"00000052",x"00000052",x"00000053",x"00000053",x"00000054",
		x"00000054",x"00000055",x"00000056",x"00000056",x"00000057",x"00000057",x"00000058",x"00000058",
		x"00000059",x"0000005a",x"0000005a",x"0000005b",x"0000005b",x"0000005c",x"0000005d",x"0000005d",
		x"0000005e",x"0000005e",x"0000005f",x"00000060",x"00000060",x"00000061",x"00000061",x"00000062",
		x"00000063",x"00000063",x"00000064",x"00000065",x"00000065",x"00000066",x"00000066",x"00000067",
		x"00000068",x"00000068",x"00000069",x"0000006a",x"0000006a",x"0000006b",x"0000006c",x"0000006c",
		x"0000006d",x"0000006e",x"0000006e",x"0000006f",x"00000070",x"00000070",x"00000071",x"00000072",
		x"00000072",x"00000073",x"00000074",x"00000074",x"00000075",x"00000076",x"00000076",x"00000077",
		x"00000078",x"00000078",x"00000079",x"0000007a",x"0000007a",x"0000007b",x"0000007c",x"0000007c",
		x"0000007d",x"0000007e",x"0000007f",x"0000007f",x"00000080",x"00000081",x"00000081",x"00000082",
		x"00000083",x"00000083",x"00000084",x"00000085",x"00000086",x"00000086",x"00000087",x"00000088",
		x"00000089",x"00000089",x"0000008a",x"0000008b",x"0000008b",x"0000008c",x"0000008d",x"0000008e",
		x"0000008e",x"0000008f",x"00000090",x"00000091",x"00000091",x"00000092",x"00000093",x"00000094",
		x"00000094",x"00000095",x"00000096",x"00000097",x"00000098",x"00000098",x"00000099",x"0000009a",
		x"0000009b",x"0000009b",x"0000009c",x"0000009d",x"0000009e",x"0000009e",x"0000009f",x"000000a0",
		x"000000a1",x"000000a2",x"000000a2",x"000000a3",x"000000a4",x"000000a5",x"000000a6",x"000000a6",
		x"000000a7",x"000000a8",x"000000a9",x"000000aa",x"000000aa",x"000000ab",x"000000ac",x"000000ad",
		x"000000ae",x"000000af",x"000000af",x"000000b0",x"000000b1",x"000000b2",x"000000b3",x"000000b4",
		x"000000b4",x"000000b5",x"000000b6",x"000000b7",x"000000b8",x"000000b9",x"000000b9",x"000000ba",
		x"000000bb",x"000000bc",x"000000bd",x"000000be",x"000000bf",x"000000bf",x"000000c0",x"000000c1",
		x"000000c2",x"000000c3",x"000000c4",x"000000c5",x"000000c5",x"000000c6",x"000000c7",x"000000c8",
		x"000000c9",x"000000ca",x"000000cb",x"000000cc",x"000000cd",x"000000cd",x"000000ce",x"000000cf",
		x"000000d0",x"000000d1",x"000000d2",x"000000d3",x"000000d4",x"000000d5",x"000000d6",x"000000d6",
		x"000000d7",x"000000d8",x"000000d9",x"000000da",x"000000db",x"000000dc",x"000000dd",x"000000de",
		x"000000df",x"000000e0",x"000000e1",x"000000e1",x"000000e2",x"000000e3",x"000000e4",x"000000e5",
		x"000000e6",x"000000e7",x"000000e8",x"000000e9",x"000000ea",x"000000eb",x"000000ec",x"000000ed",
		x"000000ee",x"000000ef",x"000000f0",x"000000f1",x"000000f2",x"000000f3",x"000000f4",x"000000f5",
		x"000000f5",x"000000f6",x"000000f7",x"000000f8",x"000000f9",x"000000fa",x"000000fb",x"000000fc",
		x"000000fd",x"000000fe",x"000000ff",x"00000100",x"00000101",x"00000102",x"00000103",x"00000104",
		x"00000105",x"00000106",x"00000107",x"00000108",x"00000109",x"0000010a",x"0000010b",x"0000010c",
		x"0000010d",x"0000010e",x"0000010f",x"00000110",x"00000111",x"00000112",x"00000114",x"00000115",
		x"00000116",x"00000117",x"00000118",x"00000119",x"0000011a",x"0000011b",x"0000011c",x"0000011d",
		x"0000011e",x"0000011f",x"00000120",x"00000121",x"00000122",x"00000123",x"00000124",x"00000125",
		x"00000126",x"00000127",x"00000128",x"0000012a",x"0000012b",x"0000012c",x"0000012d",x"0000012e",
		x"0000012f",x"00000130",x"00000131",x"00000132",x"00000133",x"00000134",x"00000135",x"00000136",
		x"00000138",x"00000139",x"0000013a",x"0000013b",x"0000013c",x"0000013d",x"0000013e",x"0000013f",
		x"00000140",x"00000141",x"00000143",x"00000144",x"00000145",x"00000146",x"00000147",x"00000148",
		x"00000149",x"0000014a",x"0000014c",x"0000014d",x"0000014e",x"0000014f",x"00000150",x"00000151",
		x"00000152",x"00000153",x"00000155",x"00000156",x"00000157",x"00000158",x"00000159",x"0000015a",
		x"0000015b",x"0000015d",x"0000015e",x"0000015f",x"00000160",x"00000161",x"00000162",x"00000164",
		x"00000165",x"00000166",x"00000167",x"00000168",x"00000169",x"0000016b",x"0000016c",x"0000016d",
		x"0000016e",x"0000016f",x"00000170",x"00000172",x"00000173",x"00000174",x"00000175",x"00000176",
		x"00000178",x"00000179",x"0000017a",x"0000017b",x"0000017c",x"0000017e",x"0000017f",x"00000180",
		x"00000181",x"00000182",x"00000184",x"00000185",x"00000186",x"00000187",x"00000188",x"0000018a",
		x"0000018b",x"0000018c",x"0000018d",x"0000018f",x"00000190",x"00000191",x"00000192",x"00000194",
		x"00000195",x"00000196",x"00000197",x"00000199",x"0000019a",x"0000019b",x"0000019c",x"0000019d",
		x"0000019f",x"000001a0",x"000001a1",x"000001a3",x"000001a4",x"000001a5",x"000001a6",x"000001a8",
		x"000001a9",x"000001aa",x"000001ab",x"000001ad",x"000001ae",x"000001af",x"000001b0",x"000001b2",
		x"000001b3",x"000001b4",x"000001b6",x"000001b7",x"000001b8",x"000001b9",x"000001bb",x"000001bc",
		x"000001bd",x"000001bf",x"000001c0",x"000001c1",x"000001c3",x"000001c4",x"000001c5",x"000001c6",
		x"000001c8",x"000001c9",x"000001ca",x"000001cc",x"000001cd",x"000001ce",x"000001d0",x"000001d1",
		x"000001d2",x"000001d4",x"000001d5",x"000001d6",x"000001d8",x"000001d9",x"000001da",x"000001dc",
		x"000001dd",x"000001de",x"000001e0",x"000001e1",x"000001e2",x"000001e4",x"000001e5",x"000001e6",
		x"000001e8",x"000001e9",x"000001ea",x"000001ec",x"000001ed",x"000001ef",x"000001f0",x"000001f1",
		x"000001f3",x"000001f4",x"000001f5",x"000001f7",x"000001f8",x"000001f9",x"000001fb",x"000001fc",
		x"000001fe",x"000001ff",x"00000200",x"00000202",x"00000203",x"00000205",x"00000206",x"00000207",
		x"00000209",x"0000020a",x"0000020c",x"0000020d",x"0000020e",x"00000210",x"00000211",x"00000213",
		x"00000214",x"00000215",x"00000217",x"00000218",x"0000021a",x"0000021b",x"0000021c",x"0000021e",
		x"0000021f",x"00000221",x"00000222",x"00000224",x"00000225",x"00000226",x"00000228",x"00000229",
		x"0000022b",x"0000022c",x"0000022e",x"0000022f",x"00000231",x"00000232",x"00000233",x"00000235",
		x"00000236",x"00000238",x"00000239",x"0000023b",x"0000023c",x"0000023e",x"0000023f",x"00000241",
		x"00000242",x"00000243",x"00000245",x"00000246",x"00000248",x"00000249",x"0000024b",x"0000024c",
		x"0000024e",x"0000024f",x"00000251",x"00000252",x"00000254",x"00000255",x"00000257",x"00000258",
		x"0000025a",x"0000025b",x"0000025d",x"0000025e",x"00000260",x"00000261",x"00000263",x"00000264",
		x"00000266",x"00000267",x"00000269",x"0000026a",x"0000026c",x"0000026d",x"0000026f",x"00000270",
		x"00000272",x"00000273",x"00000275",x"00000276",x"00000278",x"00000279",x"0000027b",x"0000027c",
		x"0000027e",x"00000280",x"00000281",x"00000283",x"00000284",x"00000286",x"00000287",x"00000289",
		x"0000028a",x"0000028c",x"0000028d",x"0000028f",x"00000291",x"00000292",x"00000294",x"00000295",
		x"00000297",x"00000298",x"0000029a",x"0000029c",x"0000029d",x"0000029f",x"000002a0",x"000002a2",
		x"000002a3",x"000002a5",x"000002a7",x"000002a8",x"000002aa",x"000002ab",x"000002ad",x"000002ae",
		x"000002b0",x"000002b2",x"000002b3",x"000002b5",x"000002b6",x"000002b8",x"000002ba",x"000002bb",
		x"000002bd",x"000002be",x"000002c0",x"000002c2",x"000002c3",x"000002c5",x"000002c6",x"000002c8",
		x"000002ca",x"000002cb",x"000002cd",x"000002cf",x"000002d0",x"000002d2",x"000002d3",x"000002d5",
		x"000002d7",x"000002d8",x"000002da",x"000002dc",x"000002dd",x"000002df",x"000002e1",x"000002e2",
		x"000002e4",x"000002e5",x"000002e7",x"000002e9",x"000002ea",x"000002ec",x"000002ee",x"000002ef",
		x"000002f1",x"000002f3",x"000002f4",x"000002f6",x"000002f8",x"000002f9",x"000002fb",x"000002fd",
		x"000002fe",x"00000300",x"00000302",x"00000303",x"00000305",x"00000307",x"00000308",x"0000030a",
		x"0000030c",x"0000030d",x"0000030f",x"00000311",x"00000313",x"00000314",x"00000316",x"00000318",
		x"00000319",x"0000031b",x"0000031d",x"0000031e",x"00000320",x"00000322",x"00000324",x"00000325",
		x"00000327",x"00000329",x"0000032a",x"0000032c",x"0000032e",x"00000330",x"00000331",x"00000333",
		x"00000335",x"00000336",x"00000338",x"0000033a",x"0000033c",x"0000033d",x"0000033f",x"00000341",
		x"00000343",x"00000344",x"00000346",x"00000348",x"0000034a",x"0000034b",x"0000034d",x"0000034f",
		x"00000350",x"00000352",x"00000354",x"00000356",x"00000358",x"00000359",x"0000035b",x"0000035d",
		x"0000035f",x"00000360",x"00000362",x"00000364",x"00000366",x"00000367",x"00000369",x"0000036b",
		x"0000036d",x"0000036f",x"00000370",x"00000372",x"00000374",x"00000376",x"00000377",x"00000379",
		x"0000037b",x"0000037d",x"0000037f",x"00000380",x"00000382",x"00000384",x"00000386",x"00000388",
		x"00000389",x"0000038b",x"0000038d",x"0000038f",x"00000391",x"00000392",x"00000394",x"00000396",
		x"00000398",x"0000039a",x"0000039b",x"0000039d",x"0000039f",x"000003a1",x"000003a3",x"000003a5",
		x"000003a6",x"000003a8",x"000003aa",x"000003ac",x"000003ae",x"000003b0",x"000003b1",x"000003b3",
		x"000003b5",x"000003b7",x"000003b9",x"000003bb",x"000003bc",x"000003be",x"000003c0",x"000003c2",
		x"000003c4",x"000003c6",x"000003c8",x"000003c9",x"000003cb",x"000003cd",x"000003cf",x"000003d1",
		x"000003d3",x"000003d5",x"000003d7",x"000003d8",x"000003da",x"000003dc",x"000003de",x"000003e0",
		x"000003e2",x"000003e4",x"000003e6",x"000003e7",x"000003e9",x"000003eb",x"000003ed",x"000003ef",
		x"000003f1",x"000003f3",x"000003f5",x"000003f7",x"000003f8",x"000003fa",x"000003fc",x"000003fe",
		x"00000400",x"00000402",x"00000404",x"00000406",x"00000408",x"0000040a",x"0000040c",x"0000040d",
		x"0000040f",x"00000411",x"00000413",x"00000415",x"00000417",x"00000419",x"0000041b",x"0000041d",
		x"0000041f",x"00000421",x"00000423",x"00000425",x"00000426",x"00000428",x"0000042a",x"0000042c",
		x"0000042e",x"00000430",x"00000432",x"00000434",x"00000436",x"00000438",x"0000043a",x"0000043c",
		x"0000043e",x"00000440",x"00000442",x"00000444",x"00000446",x"00000448",x"0000044a",x"0000044c",
		x"0000044d",x"0000044f",x"00000451",x"00000453",x"00000455",x"00000457",x"00000459",x"0000045b",
		x"0000045d",x"0000045f",x"00000461",x"00000463",x"00000465",x"00000467",x"00000469",x"0000046b",
		x"0000046d",x"0000046f",x"00000471",x"00000473",x"00000475",x"00000477",x"00000479",x"0000047b",
		x"0000047d",x"0000047f",x"00000481",x"00000483",x"00000485",x"00000487",x"00000489",x"0000048b",
		x"0000048d",x"0000048f",x"00000491",x"00000493",x"00000495",x"00000497",x"00000499",x"0000049b",
		x"0000049d",x"0000049f",x"000004a1",x"000004a4",x"000004a6",x"000004a8",x"000004aa",x"000004ac",
		x"000004ae",x"000004b0",x"000004b2",x"000004b4",x"000004b6",x"000004b8",x"000004ba",x"000004bc",
		x"000004be",x"000004c0",x"000004c2",x"000004c4",x"000004c6",x"000004c8",x"000004ca",x"000004cc",
		x"000004cf",x"000004d1",x"000004d3",x"000004d5",x"000004d7",x"000004d9",x"000004db",x"000004dd",
		x"000004df",x"000004e1",x"000004e3",x"000004e5",x"000004e7",x"000004e9",x"000004ec",x"000004ee",
		x"000004f0",x"000004f2",x"000004f4",x"000004f6",x"000004f8",x"000004fa",x"000004fc",x"000004fe",
		x"00000500",x"00000503",x"00000505",x"00000507",x"00000509",x"0000050b",x"0000050d",x"0000050f",
		x"00000511",x"00000513",x"00000516",x"00000518",x"0000051a",x"0000051c",x"0000051e",x"00000520",
		x"00000522",x"00000524",x"00000527",x"00000529",x"0000052b",x"0000052d",x"0000052f",x"00000531",
		x"00000533",x"00000535",x"00000538",x"0000053a",x"0000053c",x"0000053e",x"00000540",x"00000542",
		x"00000544",x"00000547",x"00000549",x"0000054b",x"0000054d",x"0000054f",x"00000551",x"00000553",
		x"00000556",x"00000558",x"0000055a",x"0000055c",x"0000055e",x"00000560",x"00000563",x"00000565",
		x"00000567",x"00000569",x"0000056b",x"0000056d",x"00000570",x"00000572",x"00000574",x"00000576",
		x"00000578",x"0000057b",x"0000057d",x"0000057f",x"00000581",x"00000583",x"00000585",x"00000588",
		x"0000058a",x"0000058c",x"0000058e",x"00000590",x"00000593",x"00000595",x"00000597",x"00000599",
		x"0000059b",x"0000059e",x"000005a0",x"000005a2",x"000005a4",x"000005a6",x"000005a9",x"000005ab",
		x"000005ad",x"000005af",x"000005b2",x"000005b4",x"000005b6",x"000005b8",x"000005ba",x"000005bd",
		x"000005bf",x"000005c1",x"000005c3",x"000005c6",x"000005c8",x"000005ca",x"000005cc",x"000005ce",
		x"000005d1",x"000005d3",x"000005d5",x"000005d7",x"000005da",x"000005dc",x"000005de",x"000005e0",
		x"000005e3",x"000005e5",x"000005e7",x"000005e9",x"000005ec",x"000005ee",x"000005f0",x"000005f2",
		x"000005f5",x"000005f7",x"000005f9",x"000005fb",x"000005fe",x"00000600",x"00000602",x"00000605",
		x"00000607",x"00000609",x"0000060b",x"0000060e",x"00000610",x"00000612",x"00000614",x"00000617",
		x"00000619",x"0000061b",x"0000061e",x"00000620",x"00000622",x"00000624",x"00000627",x"00000629",
		x"0000062b",x"0000062e",x"00000630",x"00000632",x"00000634",x"00000637",x"00000639",x"0000063b",
		x"0000063e",x"00000640",x"00000642",x"00000645",x"00000647",x"00000649",x"0000064b",x"0000064e",
		x"00000650",x"00000652",x"00000655",x"00000657",x"00000659",x"0000065c",x"0000065e",x"00000660",
		x"00000663",x"00000665",x"00000667",x"0000066a",x"0000066c",x"0000066e",x"00000671",x"00000673",
		x"00000675",x"00000678",x"0000067a",x"0000067c",x"0000067f",x"00000681",x"00000683",x"00000686",
		x"00000688",x"0000068a",x"0000068d",x"0000068f",x"00000691",x"00000694",x"00000696",x"00000698",
		x"0000069b",x"0000069d",x"000006a0",x"000006a2",x"000006a4",x"000006a7",x"000006a9",x"000006ab",
		x"000006ae",x"000006b0",x"000006b2",x"000006b5",x"000006b7",x"000006ba",x"000006bc",x"000006be",
		x"000006c1",x"000006c3",x"000006c5",x"000006c8",x"000006ca",x"000006cd",x"000006cf",x"000006d1",
		x"000006d4",x"000006d6",x"000006d8",x"000006db",x"000006dd",x"000006e0",x"000006e2",x"000006e4",
		x"000006e7",x"000006e9",x"000006ec",x"000006ee",x"000006f0",x"000006f3",x"000006f5",x"000006f8",
		x"000006fa",x"000006fc",x"000006ff",x"00000701",x"00000704",x"00000706",x"00000709",x"0000070b",
		x"0000070d",x"00000710",x"00000712",x"00000715",x"00000717",x"00000719",x"0000071c",x"0000071e",
		x"00000721",x"00000723",x"00000726",x"00000728",x"0000072a",x"0000072d",x"0000072f",x"00000732",
		x"00000734",x"00000737",x"00000739",x"0000073c",x"0000073e",x"00000740",x"00000743",x"00000745",
		x"00000748",x"0000074a",x"0000074d",x"0000074f",x"00000752",x"00000754",x"00000756",x"00000759",
		x"0000075b",x"0000075e",x"00000760",x"00000763",x"00000765",x"00000768",x"0000076a",x"0000076d",
		x"0000076f",x"00000772",x"00000774",x"00000776",x"00000779",x"0000077b",x"0000077e",x"00000780",
		x"00000783",x"00000785",x"00000788",x"0000078a",x"0000078d",x"0000078f",x"00000792",x"00000794",
		x"00000797",x"00000799",x"0000079c",x"0000079e",x"000007a1",x"000007a3",x"000007a6",x"000007a8",
		x"000007ab",x"000007ad",x"000007b0",x"000007b2",x"000007b5",x"000007b7",x"000007ba",x"000007bc",
		x"000007bf",x"000007c1",x"000007c4",x"000007c6",x"000007c9",x"000007cb",x"000007ce",x"000007d0",
		x"000007d3",x"000007d5",x"000007d8",x"000007da",x"000007dd",x"000007df",x"000007e2",x"000007e4",
		x"000007e7",x"000007e9",x"000007ec",x"000007ee",x"000007f1",x"000007f3",x"000007f6",x"000007f9",
		x"000007fb",x"000007fe",x"00000800",x"00000803",x"00000805",x"00000808",x"0000080a",x"0000080d",
		x"0000080f",x"00000812",x"00000814",x"00000817",x"0000081a",x"0000081c",x"0000081f",x"00000821",
		x"00000824",x"00000826",x"00000829",x"0000082b",x"0000082e",x"00000831",x"00000833",x"00000836",
		x"00000838",x"0000083b",x"0000083d",x"00000840",x"00000842",x"00000845",x"00000848",x"0000084a",
		x"0000084d",x"0000084f",x"00000852",x"00000854",x"00000857",x"0000085a",x"0000085c",x"0000085f",
		x"00000861",x"00000864",x"00000866",x"00000869",x"0000086c",x"0000086e",x"00000871",x"00000873",
		x"00000876",x"00000879",x"0000087b",x"0000087e",x"00000880",x"00000883",x"00000886",x"00000888",
		x"0000088b",x"0000088d",x"00000890",x"00000893",x"00000895",x"00000898",x"0000089a",x"0000089d",
		x"000008a0",x"000008a2",x"000008a5",x"000008a7",x"000008aa",x"000008ad",x"000008af",x"000008b2",
		x"000008b4",x"000008b7",x"000008ba",x"000008bc",x"000008bf",x"000008c2",x"000008c4",x"000008c7",
		x"000008c9",x"000008cc",x"000008cf",x"000008d1",x"000008d4",x"000008d7",x"000008d9",x"000008dc",
		x"000008de",x"000008e1",x"000008e4",x"000008e6",x"000008e9",x"000008ec",x"000008ee",x"000008f1",
		x"000008f4",x"000008f6",x"000008f9",x"000008fb",x"000008fe",x"00000901",x"00000903",x"00000906",
		x"00000909",x"0000090b",x"0000090e",x"00000911",x"00000913",x"00000916",x"00000919",x"0000091b",
		x"0000091e",x"00000921",x"00000923",x"00000926",x"00000929",x"0000092b",x"0000092e",x"00000931",
		x"00000933",x"00000936",x"00000939",x"0000093b",x"0000093e",x"00000941",x"00000943",x"00000946",
		x"00000949",x"0000094b",x"0000094e",x"00000951",x"00000953",x"00000956",x"00000959",x"0000095b",
		x"0000095e",x"00000961",x"00000963",x"00000966",x"00000969",x"0000096b",x"0000096e",x"00000971",
		x"00000973",x"00000976",x"00000979",x"0000097c",x"0000097e",x"00000981",x"00000984",x"00000986",
		x"00000989",x"0000098c",x"0000098e",x"00000991",x"00000994",x"00000997",x"00000999",x"0000099c",
		x"0000099f",x"000009a1",x"000009a4",x"000009a7",x"000009aa",x"000009ac",x"000009af",x"000009b2",
		x"000009b4",x"000009b7",x"000009ba",x"000009bd",x"000009bf",x"000009c2",x"000009c5",x"000009c7",
		x"000009ca",x"000009cd",x"000009d0",x"000009d2",x"000009d5",x"000009d8",x"000009da",x"000009dd",
		x"000009e0",x"000009e3",x"000009e5",x"000009e8",x"000009eb",x"000009ee",x"000009f0",x"000009f3",
		x"000009f6",x"000009f9",x"000009fb",x"000009fe",x"00000a01",x"00000a04",x"00000a06",x"00000a09",
		x"00000a0c",x"00000a0f",x"00000a11",x"00000a14",x"00000a17",x"00000a1a",x"00000a1c",x"00000a1f",
		x"00000a22",x"00000a25",x"00000a27",x"00000a2a",x"00000a2d",x"00000a30",x"00000a32",x"00000a35",
		x"00000a38",x"00000a3b",x"00000a3d",x"00000a40",x"00000a43",x"00000a46",x"00000a48",x"00000a4b",
		x"00000a4e",x"00000a51",x"00000a53",x"00000a56",x"00000a59",x"00000a5c",x"00000a5f",x"00000a61",
		x"00000a64",x"00000a67",x"00000a6a",x"00000a6c",x"00000a6f",x"00000a72",x"00000a75",x"00000a78",
		x"00000a7a",x"00000a7d",x"00000a80",x"00000a83",x"00000a86",x"00000a88",x"00000a8b",x"00000a8e",
		x"00000a91",x"00000a93",x"00000a96",x"00000a99",x"00000a9c",x"00000a9f",x"00000aa1",x"00000aa4",
		x"00000aa7",x"00000aaa",x"00000aad",x"00000aaf",x"00000ab2",x"00000ab5",x"00000ab8",x"00000abb",
		x"00000abd",x"00000ac0",x"00000ac3",x"00000ac6",x"00000ac9",x"00000acb",x"00000ace",x"00000ad1",
		x"00000ad4",x"00000ad7",x"00000ada",x"00000adc",x"00000adf",x"00000ae2",x"00000ae5",x"00000ae8",
		x"00000aea",x"00000aed",x"00000af0",x"00000af3",x"00000af6",x"00000af9",x"00000afb",x"00000afe",
		x"00000b01",x"00000b04",x"00000b07",x"00000b0a",x"00000b0c",x"00000b0f",x"00000b12",x"00000b15",
		x"00000b18",x"00000b1b",x"00000b1d",x"00000b20",x"00000b23",x"00000b26",x"00000b29",x"00000b2c",
		x"00000b2e",x"00000b31",x"00000b34",x"00000b37",x"00000b3a",x"00000b3d",x"00000b3f",x"00000b42",
		x"00000b45",x"00000b48",x"00000b4b",x"00000b4e",x"00000b51",x"00000b53",x"00000b56",x"00000b59",
		x"00000b5c",x"00000b5f",x"00000b62",x"00000b64",x"00000b67",x"00000b6a",x"00000b6d",x"00000b70",
		x"00000b73",x"00000b76",x"00000b79",x"00000b7b",x"00000b7e",x"00000b81",x"00000b84",x"00000b87",
		x"00000b8a",x"00000b8d",x"00000b8f",x"00000b92",x"00000b95",x"00000b98",x"00000b9b",x"00000b9e",
		x"00000ba1",x"00000ba4",x"00000ba6",x"00000ba9",x"00000bac",x"00000baf",x"00000bb2",x"00000bb5",
		x"00000bb8",x"00000bbb",x"00000bbd",x"00000bc0",x"00000bc3",x"00000bc6",x"00000bc9",x"00000bcc",
		x"00000bcf",x"00000bd2",x"00000bd5",x"00000bd7",x"00000bda",x"00000bdd",x"00000be0",x"00000be3",
		x"00000be6",x"00000be9",x"00000bec",x"00000bef",x"00000bf1",x"00000bf4",x"00000bf7",x"00000bfa",
		x"00000bfd",x"00000c00",x"00000c03",x"00000c06",x"00000c09",x"00000c0b",x"00000c0e",x"00000c11",
		x"00000c14",x"00000c17",x"00000c1a",x"00000c1d",x"00000c20",x"00000c23",x"00000c26",x"00000c29",
		x"00000c2b",x"00000c2e",x"00000c31",x"00000c34",x"00000c37",x"00000c3a",x"00000c3d",x"00000c40",
		x"00000c43",x"00000c46",x"00000c49",x"00000c4c",x"00000c4e",x"00000c51",x"00000c54",x"00000c57",
		x"00000c5a",x"00000c5d",x"00000c60",x"00000c63",x"00000c66",x"00000c69",x"00000c6c",x"00000c6f",
		x"00000c72",x"00000c74",x"00000c77",x"00000c7a",x"00000c7d",x"00000c80",x"00000c83",x"00000c86",
		x"00000c89",x"00000c8c",x"00000c8f",x"00000c92",x"00000c95",x"00000c98",x"00000c9b",x"00000c9e",
		x"00000ca0",x"00000ca3",x"00000ca6",x"00000ca9",x"00000cac",x"00000caf",x"00000cb2",x"00000cb5",
		x"00000cb8",x"00000cbb",x"00000cbe",x"00000cc1",x"00000cc4",x"00000cc7",x"00000cca",x"00000ccd",
		x"00000cd0",x"00000cd3",x"00000cd5",x"00000cd8",x"00000cdb",x"00000cde",x"00000ce1",x"00000ce4",
		x"00000ce7",x"00000cea",x"00000ced",x"00000cf0",x"00000cf3",x"00000cf6",x"00000cf9",x"00000cfc",
		x"00000cff",x"00000d02",x"00000d05",x"00000d08",x"00000d0b",x"00000d0e",x"00000d11",x"00000d14",
		x"00000d17",x"00000d1a",x"00000d1c",x"00000d1f",x"00000d22",x"00000d25",x"00000d28",x"00000d2b",
		x"00000d2e",x"00000d31",x"00000d34",x"00000d37",x"00000d3a",x"00000d3d",x"00000d40",x"00000d43",
		x"00000d46",x"00000d49",x"00000d4c",x"00000d4f",x"00000d52",x"00000d55",x"00000d58",x"00000d5b",
		x"00000d5e",x"00000d61",x"00000d64",x"00000d67",x"00000d6a",x"00000d6d",x"00000d70",x"00000d73",
		x"00000d76",x"00000d79",x"00000d7c",x"00000d7f",x"00000d82",x"00000d85",x"00000d88",x"00000d8b",
		x"00000d8e",x"00000d91",x"00000d94",x"00000d97",x"00000d9a",x"00000d9d",x"00000da0",x"00000da3",
		x"00000da6",x"00000da9",x"00000dac",x"00000daf",x"00000db2",x"00000db5",x"00000db8",x"00000dbb",
		x"00000dbe",x"00000dc1",x"00000dc4",x"00000dc7",x"00000dca",x"00000dcd",x"00000dd0",x"00000dd3",
		x"00000dd6",x"00000dd9",x"00000ddc",x"00000ddf",x"00000de2",x"00000de5",x"00000de8",x"00000deb",
		x"00000dee",x"00000df1",x"00000df4",x"00000df7",x"00000dfa",x"00000dfd",x"00000e00",x"00000e03",
		x"00000e06",x"00000e09",x"00000e0c",x"00000e0f",x"00000e12",x"00000e15",x"00000e18",x"00000e1b",
		x"00000e1e",x"00000e21",x"00000e24",x"00000e27",x"00000e2a",x"00000e2d",x"00000e30",x"00000e33",
		x"00000e36",x"00000e39",x"00000e3c",x"00000e3f",x"00000e42",x"00000e45",x"00000e48",x"00000e4b",
		x"00000e4e",x"00000e51",x"00000e54",x"00000e57",x"00000e5a",x"00000e5d",x"00000e61",x"00000e64",
		x"00000e67",x"00000e6a",x"00000e6d",x"00000e70",x"00000e73",x"00000e76",x"00000e79",x"00000e7c",
		x"00000e7f",x"00000e82",x"00000e85",x"00000e88",x"00000e8b",x"00000e8e",x"00000e91",x"00000e94",
		x"00000e97",x"00000e9a",x"00000e9d",x"00000ea0",x"00000ea3",x"00000ea6",x"00000ea9",x"00000eac",
		x"00000eaf",x"00000eb3",x"00000eb6",x"00000eb9",x"00000ebc",x"00000ebf",x"00000ec2",x"00000ec5",
		x"00000ec8",x"00000ecb",x"00000ece",x"00000ed1",x"00000ed4",x"00000ed7",x"00000eda",x"00000edd",
		x"00000ee0",x"00000ee3",x"00000ee6",x"00000ee9",x"00000eec",x"00000eef",x"00000ef3",x"00000ef6",
		x"00000ef9",x"00000efc",x"00000eff",x"00000f02",x"00000f05",x"00000f08",x"00000f0b",x"00000f0e",
		x"00000f11",x"00000f14",x"00000f17",x"00000f1a",x"00000f1d",x"00000f20",x"00000f23",x"00000f27",
		x"00000f2a",x"00000f2d",x"00000f30",x"00000f33",x"00000f36",x"00000f39",x"00000f3c",x"00000f3f",
		x"00000f42",x"00000f45",x"00000f48",x"00000f4b",x"00000f4e",x"00000f51",x"00000f55",x"00000f58",
		x"00000f5b",x"00000f5e",x"00000f61",x"00000f64",x"00000f67",x"00000f6a",x"00000f6d",x"00000f70",
		x"00000f73",x"00000f76",x"00000f79",x"00000f7c",x"00000f80",x"00000f83",x"00000f86",x"00000f89",
		x"00000f8c",x"00000f8f",x"00000f92",x"00000f95",x"00000f98",x"00000f9b",x"00000f9e",x"00000fa1",
		x"00000fa4",x"00000fa8",x"00000fab",x"00000fae",x"00000fb1",x"00000fb4",x"00000fb7",x"00000fba",
		x"00000fbd",x"00000fc0",x"00000fc3",x"00000fc6",x"00000fc9",x"00000fcc",x"00000fd0",x"00000fd3",
		x"00000fd6",x"00000fd9",x"00000fdc",x"00000fdf",x"00000fe2",x"00000fe5",x"00000fe8",x"00000feb",
		x"00000fee",x"00000ff2",x"00000ff5",x"00000ff8",x"00000ffb",x"00000ffe",x"00001001",x"00001004",
		x"00001007",x"0000100a",x"0000100d",x"00001010",x"00001014",x"00001017",x"0000101a",x"0000101d",
		x"00001020",x"00001023",x"00001026",x"00001029",x"0000102c",x"0000102f",x"00001032",x"00001036",
		x"00001039",x"0000103c",x"0000103f",x"00001042",x"00001045",x"00001048",x"0000104b",x"0000104e",
		x"00001051",x"00001055",x"00001058",x"0000105b",x"0000105e",x"00001061",x"00001064",x"00001067",
		x"0000106a",x"0000106d",x"00001070",x"00001074",x"00001077",x"0000107a",x"0000107d",x"00001080",
		x"00001083",x"00001086",x"00001089",x"0000108c",x"0000108f",x"00001093",x"00001096",x"00001099",
		x"0000109c",x"0000109f",x"000010a2",x"000010a5",x"000010a8",x"000010ab",x"000010af",x"000010b2",
		x"000010b5",x"000010b8",x"000010bb",x"000010be",x"000010c1",x"000010c4",x"000010c7",x"000010cb",
		x"000010ce",x"000010d1",x"000010d4",x"000010d7",x"000010da",x"000010dd",x"000010e0",x"000010e3",
		x"000010e7",x"000010ea",x"000010ed",x"000010f0",x"000010f3",x"000010f6",x"000010f9",x"000010fc",
		x"000010ff",x"00001103",x"00001106",x"00001109",x"0000110c",x"0000110f",x"00001112",x"00001115",
		x"00001118",x"0000111c",x"0000111f",x"00001122",x"00001125",x"00001128",x"0000112b",x"0000112e",
		x"00001131",x"00001134",x"00001138",x"0000113b",x"0000113e",x"00001141",x"00001144",x"00001147",
		x"0000114a",x"0000114d",x"00001151",x"00001154",x"00001157",x"0000115a",x"0000115d",x"00001160",
		x"00001163",x"00001166",x"0000116a",x"0000116d",x"00001170",x"00001173",x"00001176",x"00001179",
		x"0000117c",x"0000117f",x"00001183",x"00001186",x"00001189",x"0000118c",x"0000118f",x"00001192",
		x"00001195",x"00001198",x"0000119c",x"0000119f",x"000011a2",x"000011a5",x"000011a8",x"000011ab",
		x"000011ae",x"000011b1",x"000011b5",x"000011b8",x"000011bb",x"000011be",x"000011c1",x"000011c4",
		x"000011c7",x"000011ca",x"000011ce",x"000011d1",x"000011d4",x"000011d7",x"000011da",x"000011dd",
		x"000011e0",x"000011e3",x"000011e7",x"000011ea",x"000011ed",x"000011f0",x"000011f3",x"000011f6",
		x"000011f9",x"000011fd",x"00001200",x"00001203",x"00001206",x"00001209",x"0000120c",x"0000120f",
		x"00001212",x"00001216",x"00001219",x"0000121c",x"0000121f",x"00001222",x"00001225",x"00001228",
		x"0000122c",x"0000122f",x"00001232",x"00001235",x"00001238",x"0000123b",x"0000123e",x"00001241",
		x"00001245",x"00001248",x"0000124b",x"0000124e",x"00001251",x"00001254",x"00001257",x"0000125b",
		x"0000125e",x"00001261",x"00001264",x"00001267",x"0000126a",x"0000126d",x"00001271",x"00001274",
		x"00001277",x"0000127a",x"0000127d",x"00001280",x"00001283",x"00001286",x"0000128a",x"0000128d",
		x"00001290",x"00001293",x"00001296",x"00001299",x"0000129c",x"000012a0",x"000012a3",x"000012a6",
		x"000012a9",x"000012ac",x"000012af",x"000012b2",x"000012b6",x"000012b9",x"000012bc",x"000012bf",
		x"000012c2",x"000012c5",x"000012c8",x"000012cc",x"000012cf",x"000012d2",x"000012d5",x"000012d8",
		x"000012db",x"000012de",x"000012e2",x"000012e5",x"000012e8",x"000012eb",x"000012ee",x"000012f1",
		x"000012f4",x"000012f7",x"000012fb",x"000012fe",x"00001301",x"00001304",x"00001307",x"0000130a",
		x"0000130d",x"00001311",x"00001314",x"00001317",x"0000131a",x"0000131d",x"00001320",x"00001323",
		x"00001327",x"0000132a",x"0000132d",x"00001330",x"00001333",x"00001336",x"00001339",x"0000133d",
		x"00001340",x"00001343",x"00001346",x"00001349",x"0000134c",x"0000134f",x"00001353",x"00001356",
		x"00001359",x"0000135c",x"0000135f",x"00001362",x"00001365",x"00001369",x"0000136c",x"0000136f",
		x"00001372",x"00001375",x"00001378",x"0000137b",x"0000137f",x"00001382",x"00001385",x"00001388"
	);
	

begin
    
	process (clk)
		variable counter:	std_logic_vector(32-1 downto 0) := (others => '0');
		variable index: natural := 1;
		variable cociente : natural :=1;
		variable resto : integer :=0;
	begin
		if (rising_edge(clk)) then
			counter := counter + 10000;--Lo cambio a 200 para 20ns

			if (counter >= frq) then
				cociente:=((to_integer(unsigned(std_logic_vector(counter))))/(to_integer(unsigned(std_logic_vector(frq)))));
				index:=index + cociente;
				resto:=((to_integer(unsigned(std_logic_vector(counter))))rem(to_integer(unsigned(std_logic_vector(frq)))));
				counter:= std_logic_vector(to_unsigned(resto, 32));
				--counter := (others => '0');
			end if;

			-- if index > 100 reset it to 1
			if (index > 10000) then
				index := 1;
			end if;
		end if;
		pwm_ctrl <= data(index);
	end process;

end Behavioral;